VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO DAC
  CLASS BLOCK ;
  FOREIGN DAC ;
  ORIGIN 12.310 12.870 ;
  SIZE 58.055 BY 28.630 ;
  PIN D3
    ANTENNAGATEAREA 1.080000 ;
    PORT
      LAYER met1 ;
        RECT 29.570 10.060 30.570 11.060 ;
    END
  END D3
  PIN D2
    ANTENNAGATEAREA 1.080000 ;
    PORT
      LAYER met1 ;
        RECT 23.090 9.860 24.090 10.860 ;
    END
  END D2
  PIN D0
    ANTENNAGATEAREA 1.080000 ;
    PORT
      LAYER met1 ;
        RECT 10.440 10.620 11.440 11.620 ;
    END
  END D0
  PIN D1
    ANTENNAGATEAREA 1.080000 ;
    PORT
      LAYER met1 ;
        RECT 16.670 10.220 17.670 11.220 ;
    END
  END D1
  PIN Vref
    PORT
      LAYER met1 ;
        RECT -12.310 -4.710 -11.310 -3.710 ;
    END
  END Vref
  PIN OUT
    ANTENNADIFFAREA 4.760000 ;
    PORT
      LAYER met1 ;
        RECT 32.060 9.180 33.060 10.180 ;
    END
  END OUT
  PIN VDD
    PORT
      LAYER met1 ;
        RECT 44.745 8.375 45.745 9.375 ;
    END
  END VDD
  PIN VSS
    ANTENNADIFFAREA 64.836502 ;
    PORT
      LAYER met1 ;
        RECT 13.710 -12.870 14.850 -11.490 ;
    END
  END VSS
  OBS
      LAYER nwell ;
        RECT -9.700 -8.600 41.410 15.760 ;
      LAYER li1 ;
        RECT -9.520 -8.600 41.230 15.580 ;
      LAYER met1 ;
        RECT -11.310 11.900 44.745 14.900 ;
        RECT -11.310 10.340 10.160 11.900 ;
        RECT 11.720 11.500 44.745 11.900 ;
        RECT 11.720 10.340 16.390 11.500 ;
        RECT -11.310 9.940 16.390 10.340 ;
        RECT 17.950 11.340 44.745 11.500 ;
        RECT 17.950 11.140 29.290 11.340 ;
        RECT 17.950 9.940 22.810 11.140 ;
        RECT -11.310 9.580 22.810 9.940 ;
        RECT 24.370 9.780 29.290 11.140 ;
        RECT 30.850 10.460 44.745 11.340 ;
        RECT 30.850 9.780 31.780 10.460 ;
        RECT 24.370 9.580 31.780 9.780 ;
        RECT -11.310 8.900 31.780 9.580 ;
        RECT 33.340 9.655 44.745 10.460 ;
        RECT 33.340 8.900 44.465 9.655 ;
        RECT -11.310 8.095 44.465 8.900 ;
        RECT -11.310 -3.430 44.745 8.095 ;
        RECT -11.030 -4.990 44.745 -3.430 ;
        RECT -11.310 -11.210 44.745 -4.990 ;
        RECT -11.310 -11.490 13.430 -11.210 ;
        RECT 15.130 -11.490 44.745 -11.210 ;
      LAYER met2 ;
        RECT -0.520 -7.660 42.150 10.280 ;
  END
END DAC
END LIBRARY

