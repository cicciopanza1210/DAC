magic
tech sky130A
magscale 1 2
timestamp 1751989567
<< error_p >>
rect -1037 360 -979 366
rect -845 360 -787 366
rect -653 360 -595 366
rect -461 360 -403 366
rect -269 360 -211 366
rect -77 360 -19 366
rect 115 360 173 366
rect 307 360 365 366
rect 499 360 557 366
rect 691 360 749 366
rect 883 360 941 366
rect 1075 360 1133 366
rect -1037 326 -1025 360
rect -845 326 -833 360
rect -653 326 -641 360
rect -461 326 -449 360
rect -269 326 -257 360
rect -77 326 -65 360
rect 115 326 127 360
rect 307 326 319 360
rect 499 326 511 360
rect 691 326 703 360
rect 883 326 895 360
rect 1075 326 1087 360
rect -1037 320 -979 326
rect -845 320 -787 326
rect -653 320 -595 326
rect -461 320 -403 326
rect -269 320 -211 326
rect -77 320 -19 326
rect 115 320 173 326
rect 307 320 365 326
rect 499 320 557 326
rect 691 320 749 326
rect 883 320 941 326
rect 1075 320 1133 326
rect -1133 -326 -1075 -320
rect -941 -326 -883 -320
rect -749 -326 -691 -320
rect -557 -326 -499 -320
rect -365 -326 -307 -320
rect -173 -326 -115 -320
rect 19 -326 77 -320
rect 211 -326 269 -320
rect 403 -326 461 -320
rect 595 -326 653 -320
rect 787 -326 845 -320
rect 979 -326 1037 -320
rect -1133 -360 -1121 -326
rect -941 -360 -929 -326
rect -749 -360 -737 -326
rect -557 -360 -545 -326
rect -365 -360 -353 -326
rect -173 -360 -161 -326
rect 19 -360 31 -326
rect 211 -360 223 -326
rect 403 -360 415 -326
rect 595 -360 607 -326
rect 787 -360 799 -326
rect 979 -360 991 -326
rect -1133 -366 -1075 -360
rect -941 -366 -883 -360
rect -749 -366 -691 -360
rect -557 -366 -499 -360
rect -365 -366 -307 -360
rect -173 -366 -115 -360
rect 19 -366 77 -360
rect 211 -366 269 -360
rect 403 -366 461 -360
rect 595 -366 653 -360
rect 787 -366 845 -360
rect 979 -366 1037 -360
<< pwell >>
rect -1319 -498 1319 498
<< nmoslvt >>
rect -1122 -288 -1086 288
rect -1026 -288 -990 288
rect -930 -288 -894 288
rect -834 -288 -798 288
rect -738 -288 -702 288
rect -642 -288 -606 288
rect -546 -288 -510 288
rect -450 -288 -414 288
rect -354 -288 -318 288
rect -258 -288 -222 288
rect -162 -288 -126 288
rect -66 -288 -30 288
rect 30 -288 66 288
rect 126 -288 162 288
rect 222 -288 258 288
rect 318 -288 354 288
rect 414 -288 450 288
rect 510 -288 546 288
rect 606 -288 642 288
rect 702 -288 738 288
rect 798 -288 834 288
rect 894 -288 930 288
rect 990 -288 1026 288
rect 1086 -288 1122 288
<< ndiff >>
rect -1181 276 -1122 288
rect -1181 -276 -1169 276
rect -1135 -276 -1122 276
rect -1181 -288 -1122 -276
rect -1086 276 -1026 288
rect -1086 -276 -1073 276
rect -1039 -276 -1026 276
rect -1086 -288 -1026 -276
rect -990 276 -930 288
rect -990 -276 -977 276
rect -943 -276 -930 276
rect -990 -288 -930 -276
rect -894 276 -834 288
rect -894 -276 -881 276
rect -847 -276 -834 276
rect -894 -288 -834 -276
rect -798 276 -738 288
rect -798 -276 -785 276
rect -751 -276 -738 276
rect -798 -288 -738 -276
rect -702 276 -642 288
rect -702 -276 -689 276
rect -655 -276 -642 276
rect -702 -288 -642 -276
rect -606 276 -546 288
rect -606 -276 -593 276
rect -559 -276 -546 276
rect -606 -288 -546 -276
rect -510 276 -450 288
rect -510 -276 -497 276
rect -463 -276 -450 276
rect -510 -288 -450 -276
rect -414 276 -354 288
rect -414 -276 -401 276
rect -367 -276 -354 276
rect -414 -288 -354 -276
rect -318 276 -258 288
rect -318 -276 -305 276
rect -271 -276 -258 276
rect -318 -288 -258 -276
rect -222 276 -162 288
rect -222 -276 -209 276
rect -175 -276 -162 276
rect -222 -288 -162 -276
rect -126 276 -66 288
rect -126 -276 -113 276
rect -79 -276 -66 276
rect -126 -288 -66 -276
rect -30 276 30 288
rect -30 -276 -17 276
rect 17 -276 30 276
rect -30 -288 30 -276
rect 66 276 126 288
rect 66 -276 79 276
rect 113 -276 126 276
rect 66 -288 126 -276
rect 162 276 222 288
rect 162 -276 175 276
rect 209 -276 222 276
rect 162 -288 222 -276
rect 258 276 318 288
rect 258 -276 271 276
rect 305 -276 318 276
rect 258 -288 318 -276
rect 354 276 414 288
rect 354 -276 367 276
rect 401 -276 414 276
rect 354 -288 414 -276
rect 450 276 510 288
rect 450 -276 463 276
rect 497 -276 510 276
rect 450 -288 510 -276
rect 546 276 606 288
rect 546 -276 559 276
rect 593 -276 606 276
rect 546 -288 606 -276
rect 642 276 702 288
rect 642 -276 655 276
rect 689 -276 702 276
rect 642 -288 702 -276
rect 738 276 798 288
rect 738 -276 751 276
rect 785 -276 798 276
rect 738 -288 798 -276
rect 834 276 894 288
rect 834 -276 847 276
rect 881 -276 894 276
rect 834 -288 894 -276
rect 930 276 990 288
rect 930 -276 943 276
rect 977 -276 990 276
rect 930 -288 990 -276
rect 1026 276 1086 288
rect 1026 -276 1039 276
rect 1073 -276 1086 276
rect 1026 -288 1086 -276
rect 1122 276 1181 288
rect 1122 -276 1135 276
rect 1169 -276 1181 276
rect 1122 -288 1181 -276
<< ndiffc >>
rect -1169 -276 -1135 276
rect -1073 -276 -1039 276
rect -977 -276 -943 276
rect -881 -276 -847 276
rect -785 -276 -751 276
rect -689 -276 -655 276
rect -593 -276 -559 276
rect -497 -276 -463 276
rect -401 -276 -367 276
rect -305 -276 -271 276
rect -209 -276 -175 276
rect -113 -276 -79 276
rect -17 -276 17 276
rect 79 -276 113 276
rect 175 -276 209 276
rect 271 -276 305 276
rect 367 -276 401 276
rect 463 -276 497 276
rect 559 -276 593 276
rect 655 -276 689 276
rect 751 -276 785 276
rect 847 -276 881 276
rect 943 -276 977 276
rect 1039 -276 1073 276
rect 1135 -276 1169 276
<< psubdiff >>
rect -1283 428 -1187 462
rect 1187 428 1283 462
rect -1283 366 -1249 428
rect 1249 366 1283 428
rect -1283 -428 -1249 -366
rect 1249 -428 1283 -366
rect -1283 -462 -1187 -428
rect 1187 -462 1283 -428
<< psubdiffcont >>
rect -1187 428 1187 462
rect -1283 -366 -1249 366
rect 1249 -366 1283 366
rect -1187 -462 1187 -428
<< poly >>
rect -1041 360 -975 376
rect -1041 326 -1025 360
rect -991 326 -975 360
rect -1122 288 -1086 314
rect -1041 310 -975 326
rect -849 360 -783 376
rect -849 326 -833 360
rect -799 326 -783 360
rect -1026 288 -990 310
rect -930 288 -894 314
rect -849 310 -783 326
rect -657 360 -591 376
rect -657 326 -641 360
rect -607 326 -591 360
rect -834 288 -798 310
rect -738 288 -702 314
rect -657 310 -591 326
rect -465 360 -399 376
rect -465 326 -449 360
rect -415 326 -399 360
rect -642 288 -606 310
rect -546 288 -510 314
rect -465 310 -399 326
rect -273 360 -207 376
rect -273 326 -257 360
rect -223 326 -207 360
rect -450 288 -414 310
rect -354 288 -318 314
rect -273 310 -207 326
rect -81 360 -15 376
rect -81 326 -65 360
rect -31 326 -15 360
rect -258 288 -222 310
rect -162 288 -126 314
rect -81 310 -15 326
rect 111 360 177 376
rect 111 326 127 360
rect 161 326 177 360
rect -66 288 -30 310
rect 30 288 66 314
rect 111 310 177 326
rect 303 360 369 376
rect 303 326 319 360
rect 353 326 369 360
rect 126 288 162 310
rect 222 288 258 314
rect 303 310 369 326
rect 495 360 561 376
rect 495 326 511 360
rect 545 326 561 360
rect 318 288 354 310
rect 414 288 450 314
rect 495 310 561 326
rect 687 360 753 376
rect 687 326 703 360
rect 737 326 753 360
rect 510 288 546 310
rect 606 288 642 314
rect 687 310 753 326
rect 879 360 945 376
rect 879 326 895 360
rect 929 326 945 360
rect 702 288 738 310
rect 798 288 834 314
rect 879 310 945 326
rect 1071 360 1137 376
rect 1071 326 1087 360
rect 1121 326 1137 360
rect 894 288 930 310
rect 990 288 1026 314
rect 1071 310 1137 326
rect 1086 288 1122 310
rect -1122 -310 -1086 -288
rect -1137 -326 -1071 -310
rect -1026 -314 -990 -288
rect -930 -310 -894 -288
rect -1137 -360 -1121 -326
rect -1087 -360 -1071 -326
rect -1137 -376 -1071 -360
rect -945 -326 -879 -310
rect -834 -314 -798 -288
rect -738 -310 -702 -288
rect -945 -360 -929 -326
rect -895 -360 -879 -326
rect -945 -376 -879 -360
rect -753 -326 -687 -310
rect -642 -314 -606 -288
rect -546 -310 -510 -288
rect -753 -360 -737 -326
rect -703 -360 -687 -326
rect -753 -376 -687 -360
rect -561 -326 -495 -310
rect -450 -314 -414 -288
rect -354 -310 -318 -288
rect -561 -360 -545 -326
rect -511 -360 -495 -326
rect -561 -376 -495 -360
rect -369 -326 -303 -310
rect -258 -314 -222 -288
rect -162 -310 -126 -288
rect -369 -360 -353 -326
rect -319 -360 -303 -326
rect -369 -376 -303 -360
rect -177 -326 -111 -310
rect -66 -314 -30 -288
rect 30 -310 66 -288
rect -177 -360 -161 -326
rect -127 -360 -111 -326
rect -177 -376 -111 -360
rect 15 -326 81 -310
rect 126 -314 162 -288
rect 222 -310 258 -288
rect 15 -360 31 -326
rect 65 -360 81 -326
rect 15 -376 81 -360
rect 207 -326 273 -310
rect 318 -314 354 -288
rect 414 -310 450 -288
rect 207 -360 223 -326
rect 257 -360 273 -326
rect 207 -376 273 -360
rect 399 -326 465 -310
rect 510 -314 546 -288
rect 606 -310 642 -288
rect 399 -360 415 -326
rect 449 -360 465 -326
rect 399 -376 465 -360
rect 591 -326 657 -310
rect 702 -314 738 -288
rect 798 -310 834 -288
rect 591 -360 607 -326
rect 641 -360 657 -326
rect 591 -376 657 -360
rect 783 -326 849 -310
rect 894 -314 930 -288
rect 990 -310 1026 -288
rect 783 -360 799 -326
rect 833 -360 849 -326
rect 783 -376 849 -360
rect 975 -326 1041 -310
rect 1086 -314 1122 -288
rect 975 -360 991 -326
rect 1025 -360 1041 -326
rect 975 -376 1041 -360
<< polycont >>
rect -1025 326 -991 360
rect -833 326 -799 360
rect -641 326 -607 360
rect -449 326 -415 360
rect -257 326 -223 360
rect -65 326 -31 360
rect 127 326 161 360
rect 319 326 353 360
rect 511 326 545 360
rect 703 326 737 360
rect 895 326 929 360
rect 1087 326 1121 360
rect -1121 -360 -1087 -326
rect -929 -360 -895 -326
rect -737 -360 -703 -326
rect -545 -360 -511 -326
rect -353 -360 -319 -326
rect -161 -360 -127 -326
rect 31 -360 65 -326
rect 223 -360 257 -326
rect 415 -360 449 -326
rect 607 -360 641 -326
rect 799 -360 833 -326
rect 991 -360 1025 -326
<< locali >>
rect -1283 428 -1187 462
rect 1187 428 1283 462
rect -1283 366 -1249 428
rect 1249 366 1283 428
rect -1041 326 -1025 360
rect -991 326 -975 360
rect -849 326 -833 360
rect -799 326 -783 360
rect -657 326 -641 360
rect -607 326 -591 360
rect -465 326 -449 360
rect -415 326 -399 360
rect -273 326 -257 360
rect -223 326 -207 360
rect -81 326 -65 360
rect -31 326 -15 360
rect 111 326 127 360
rect 161 326 177 360
rect 303 326 319 360
rect 353 326 369 360
rect 495 326 511 360
rect 545 326 561 360
rect 687 326 703 360
rect 737 326 753 360
rect 879 326 895 360
rect 929 326 945 360
rect 1071 326 1087 360
rect 1121 326 1137 360
rect -1169 276 -1135 292
rect -1169 -292 -1135 -276
rect -1073 276 -1039 292
rect -1073 -292 -1039 -276
rect -977 276 -943 292
rect -977 -292 -943 -276
rect -881 276 -847 292
rect -881 -292 -847 -276
rect -785 276 -751 292
rect -785 -292 -751 -276
rect -689 276 -655 292
rect -689 -292 -655 -276
rect -593 276 -559 292
rect -593 -292 -559 -276
rect -497 276 -463 292
rect -497 -292 -463 -276
rect -401 276 -367 292
rect -401 -292 -367 -276
rect -305 276 -271 292
rect -305 -292 -271 -276
rect -209 276 -175 292
rect -209 -292 -175 -276
rect -113 276 -79 292
rect -113 -292 -79 -276
rect -17 276 17 292
rect -17 -292 17 -276
rect 79 276 113 292
rect 79 -292 113 -276
rect 175 276 209 292
rect 175 -292 209 -276
rect 271 276 305 292
rect 271 -292 305 -276
rect 367 276 401 292
rect 367 -292 401 -276
rect 463 276 497 292
rect 463 -292 497 -276
rect 559 276 593 292
rect 559 -292 593 -276
rect 655 276 689 292
rect 655 -292 689 -276
rect 751 276 785 292
rect 751 -292 785 -276
rect 847 276 881 292
rect 847 -292 881 -276
rect 943 276 977 292
rect 943 -292 977 -276
rect 1039 276 1073 292
rect 1039 -292 1073 -276
rect 1135 276 1169 292
rect 1135 -292 1169 -276
rect -1137 -360 -1121 -326
rect -1087 -360 -1071 -326
rect -945 -360 -929 -326
rect -895 -360 -879 -326
rect -753 -360 -737 -326
rect -703 -360 -687 -326
rect -561 -360 -545 -326
rect -511 -360 -495 -326
rect -369 -360 -353 -326
rect -319 -360 -303 -326
rect -177 -360 -161 -326
rect -127 -360 -111 -326
rect 15 -360 31 -326
rect 65 -360 81 -326
rect 207 -360 223 -326
rect 257 -360 273 -326
rect 399 -360 415 -326
rect 449 -360 465 -326
rect 591 -360 607 -326
rect 641 -360 657 -326
rect 783 -360 799 -326
rect 833 -360 849 -326
rect 975 -360 991 -326
rect 1025 -360 1041 -326
rect -1283 -428 -1249 -366
rect 1249 -428 1283 -366
rect -1283 -462 -1187 -428
rect 1187 -462 1283 -428
<< viali >>
rect -1025 326 -991 360
rect -833 326 -799 360
rect -641 326 -607 360
rect -449 326 -415 360
rect -257 326 -223 360
rect -65 326 -31 360
rect 127 326 161 360
rect 319 326 353 360
rect 511 326 545 360
rect 703 326 737 360
rect 895 326 929 360
rect 1087 326 1121 360
rect -1169 -276 -1135 276
rect -1073 -276 -1039 276
rect -977 -276 -943 276
rect -881 -276 -847 276
rect -785 -276 -751 276
rect -689 -276 -655 276
rect -593 -276 -559 276
rect -497 -276 -463 276
rect -401 -276 -367 276
rect -305 -276 -271 276
rect -209 -276 -175 276
rect -113 -276 -79 276
rect -17 -276 17 276
rect 79 -276 113 276
rect 175 -276 209 276
rect 271 -276 305 276
rect 367 -276 401 276
rect 463 -276 497 276
rect 559 -276 593 276
rect 655 -276 689 276
rect 751 -276 785 276
rect 847 -276 881 276
rect 943 -276 977 276
rect 1039 -276 1073 276
rect 1135 -276 1169 276
rect -1121 -360 -1087 -326
rect -929 -360 -895 -326
rect -737 -360 -703 -326
rect -545 -360 -511 -326
rect -353 -360 -319 -326
rect -161 -360 -127 -326
rect 31 -360 65 -326
rect 223 -360 257 -326
rect 415 -360 449 -326
rect 607 -360 641 -326
rect 799 -360 833 -326
rect 991 -360 1025 -326
<< metal1 >>
rect -1037 360 -979 366
rect -1037 326 -1025 360
rect -991 326 -979 360
rect -1037 320 -979 326
rect -845 360 -787 366
rect -845 326 -833 360
rect -799 326 -787 360
rect -845 320 -787 326
rect -653 360 -595 366
rect -653 326 -641 360
rect -607 326 -595 360
rect -653 320 -595 326
rect -461 360 -403 366
rect -461 326 -449 360
rect -415 326 -403 360
rect -461 320 -403 326
rect -269 360 -211 366
rect -269 326 -257 360
rect -223 326 -211 360
rect -269 320 -211 326
rect -77 360 -19 366
rect -77 326 -65 360
rect -31 326 -19 360
rect -77 320 -19 326
rect 115 360 173 366
rect 115 326 127 360
rect 161 326 173 360
rect 115 320 173 326
rect 307 360 365 366
rect 307 326 319 360
rect 353 326 365 360
rect 307 320 365 326
rect 499 360 557 366
rect 499 326 511 360
rect 545 326 557 360
rect 499 320 557 326
rect 691 360 749 366
rect 691 326 703 360
rect 737 326 749 360
rect 691 320 749 326
rect 883 360 941 366
rect 883 326 895 360
rect 929 326 941 360
rect 883 320 941 326
rect 1075 360 1133 366
rect 1075 326 1087 360
rect 1121 326 1133 360
rect 1075 320 1133 326
rect -1175 276 -1129 288
rect -1175 -276 -1169 276
rect -1135 -276 -1129 276
rect -1175 -288 -1129 -276
rect -1079 276 -1033 288
rect -1079 -276 -1073 276
rect -1039 -276 -1033 276
rect -1079 -288 -1033 -276
rect -983 276 -937 288
rect -983 -276 -977 276
rect -943 -276 -937 276
rect -983 -288 -937 -276
rect -887 276 -841 288
rect -887 -276 -881 276
rect -847 -276 -841 276
rect -887 -288 -841 -276
rect -791 276 -745 288
rect -791 -276 -785 276
rect -751 -276 -745 276
rect -791 -288 -745 -276
rect -695 276 -649 288
rect -695 -276 -689 276
rect -655 -276 -649 276
rect -695 -288 -649 -276
rect -599 276 -553 288
rect -599 -276 -593 276
rect -559 -276 -553 276
rect -599 -288 -553 -276
rect -503 276 -457 288
rect -503 -276 -497 276
rect -463 -276 -457 276
rect -503 -288 -457 -276
rect -407 276 -361 288
rect -407 -276 -401 276
rect -367 -276 -361 276
rect -407 -288 -361 -276
rect -311 276 -265 288
rect -311 -276 -305 276
rect -271 -276 -265 276
rect -311 -288 -265 -276
rect -215 276 -169 288
rect -215 -276 -209 276
rect -175 -276 -169 276
rect -215 -288 -169 -276
rect -119 276 -73 288
rect -119 -276 -113 276
rect -79 -276 -73 276
rect -119 -288 -73 -276
rect -23 276 23 288
rect -23 -276 -17 276
rect 17 -276 23 276
rect -23 -288 23 -276
rect 73 276 119 288
rect 73 -276 79 276
rect 113 -276 119 276
rect 73 -288 119 -276
rect 169 276 215 288
rect 169 -276 175 276
rect 209 -276 215 276
rect 169 -288 215 -276
rect 265 276 311 288
rect 265 -276 271 276
rect 305 -276 311 276
rect 265 -288 311 -276
rect 361 276 407 288
rect 361 -276 367 276
rect 401 -276 407 276
rect 361 -288 407 -276
rect 457 276 503 288
rect 457 -276 463 276
rect 497 -276 503 276
rect 457 -288 503 -276
rect 553 276 599 288
rect 553 -276 559 276
rect 593 -276 599 276
rect 553 -288 599 -276
rect 649 276 695 288
rect 649 -276 655 276
rect 689 -276 695 276
rect 649 -288 695 -276
rect 745 276 791 288
rect 745 -276 751 276
rect 785 -276 791 276
rect 745 -288 791 -276
rect 841 276 887 288
rect 841 -276 847 276
rect 881 -276 887 276
rect 841 -288 887 -276
rect 937 276 983 288
rect 937 -276 943 276
rect 977 -276 983 276
rect 937 -288 983 -276
rect 1033 276 1079 288
rect 1033 -276 1039 276
rect 1073 -276 1079 276
rect 1033 -288 1079 -276
rect 1129 276 1175 288
rect 1129 -276 1135 276
rect 1169 -276 1175 276
rect 1129 -288 1175 -276
rect -1133 -326 -1075 -320
rect -1133 -360 -1121 -326
rect -1087 -360 -1075 -326
rect -1133 -366 -1075 -360
rect -941 -326 -883 -320
rect -941 -360 -929 -326
rect -895 -360 -883 -326
rect -941 -366 -883 -360
rect -749 -326 -691 -320
rect -749 -360 -737 -326
rect -703 -360 -691 -326
rect -749 -366 -691 -360
rect -557 -326 -499 -320
rect -557 -360 -545 -326
rect -511 -360 -499 -326
rect -557 -366 -499 -360
rect -365 -326 -307 -320
rect -365 -360 -353 -326
rect -319 -360 -307 -326
rect -365 -366 -307 -360
rect -173 -326 -115 -320
rect -173 -360 -161 -326
rect -127 -360 -115 -326
rect -173 -366 -115 -360
rect 19 -326 77 -320
rect 19 -360 31 -326
rect 65 -360 77 -326
rect 19 -366 77 -360
rect 211 -326 269 -320
rect 211 -360 223 -326
rect 257 -360 269 -326
rect 211 -366 269 -360
rect 403 -326 461 -320
rect 403 -360 415 -326
rect 449 -360 461 -326
rect 403 -366 461 -360
rect 595 -326 653 -320
rect 595 -360 607 -326
rect 641 -360 653 -326
rect 595 -366 653 -360
rect 787 -326 845 -320
rect 787 -360 799 -326
rect 833 -360 845 -326
rect 787 -366 845 -360
rect 979 -326 1037 -320
rect 979 -360 991 -326
rect 1025 -360 1037 -326
rect 979 -366 1037 -360
<< properties >>
string FIXED_BBOX -1266 -445 1266 445
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2.875 l 0.18 m 1 nf 24 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
