magic
tech sky130A
magscale 1 2
timestamp 1752588718
<< error_p >>
rect 7449 5454 7811 5460
rect 7449 5226 7455 5454
rect 7805 5226 7811 5454
rect 7449 5220 7811 5226
rect 5536 4225 5571 4259
rect 5537 4206 5571 4225
rect -1964 1105 -1929 1139
rect -1963 1086 -1929 1105
rect -2233 1037 -2175 1043
rect -2233 1003 -2221 1037
rect -2233 997 -2175 1003
rect -2329 527 -2271 533
rect -2137 527 -2079 533
rect -2329 493 -2317 527
rect -2137 493 -2125 527
rect -2329 487 -2271 493
rect -2137 487 -2079 493
rect -1944 391 -1929 1086
rect -1910 1052 -1875 1086
rect -1395 1052 -1360 1086
rect -1910 391 -1876 1052
rect -1394 1033 -1360 1052
rect -772 1080 -737 1087
rect -257 1080 -222 1114
rect -1664 984 -1606 990
rect -1664 950 -1652 984
rect -1664 944 -1606 950
rect -1760 474 -1702 480
rect -1568 474 -1510 480
rect -1760 440 -1748 474
rect -1568 440 -1556 474
rect -1760 434 -1702 440
rect -1568 434 -1510 440
rect -1910 357 -1895 391
rect -1375 338 -1360 1033
rect -1341 999 -1306 1033
rect -1341 338 -1307 999
rect -1095 931 -1037 937
rect -1095 897 -1083 931
rect -1095 891 -1037 897
rect -1191 421 -1133 427
rect -999 421 -941 427
rect -1191 387 -1179 421
rect -999 387 -987 421
rect -1191 381 -1133 387
rect -999 381 -941 387
rect -1341 304 -1326 338
rect -806 285 -791 1033
rect -772 285 -738 1080
rect -256 1061 -222 1080
rect -526 1012 -468 1018
rect -526 978 -514 1012
rect -526 972 -468 978
rect -622 368 -564 374
rect -430 368 -372 374
rect -622 334 -610 368
rect -430 334 -418 368
rect -622 328 -564 334
rect -430 328 -372 334
rect -772 251 -757 285
rect -237 232 -222 1061
rect -203 1027 -168 1061
rect 600 1027 635 1061
rect -203 232 -169 1027
rect 601 1024 635 1027
rect 43 959 101 965
rect 235 959 293 965
rect 427 959 485 965
rect 43 925 55 959
rect 235 925 247 959
rect 427 925 439 959
rect 43 919 101 925
rect 235 919 293 925
rect 427 919 485 925
rect -53 315 5 321
rect 139 315 197 321
rect 331 315 389 321
rect -53 281 -41 315
rect 139 281 151 315
rect 331 281 343 315
rect -53 275 5 281
rect 139 275 197 281
rect 331 275 389 281
rect -203 198 -188 232
rect 620 179 635 1024
rect 654 990 689 1024
rect 2033 997 2068 1024
rect 654 179 688 990
rect 900 922 958 928
rect 1092 922 1150 928
rect 1284 922 1342 928
rect 1476 922 1534 928
rect 1668 922 1726 928
rect 1860 922 1918 928
rect 900 888 912 922
rect 1092 888 1104 922
rect 1284 888 1296 922
rect 1476 888 1488 922
rect 1668 888 1680 922
rect 1860 888 1872 922
rect 900 882 958 888
rect 1092 882 1150 888
rect 1284 882 1342 888
rect 1476 882 1534 888
rect 1668 882 1726 888
rect 1860 882 1918 888
rect 804 262 862 268
rect 996 262 1054 268
rect 1188 262 1246 268
rect 1380 262 1438 268
rect 1572 262 1630 268
rect 1764 262 1822 268
rect 804 228 816 262
rect 996 228 1008 262
rect 1188 228 1200 262
rect 1380 228 1392 262
rect 1572 228 1584 262
rect 1764 228 1776 262
rect 804 222 862 228
rect 996 222 1054 228
rect 1188 222 1246 228
rect 1380 222 1438 228
rect 1572 222 1630 228
rect 1764 222 1822 228
rect 654 145 669 179
rect 2053 126 2068 997
rect 2087 963 2122 997
rect 2087 126 2121 963
rect 4619 902 4653 956
rect 2333 895 2391 901
rect 2525 895 2583 901
rect 2717 895 2775 901
rect 2909 895 2967 901
rect 3101 895 3159 901
rect 3293 895 3351 901
rect 3485 895 3543 901
rect 3677 895 3735 901
rect 3869 895 3927 901
rect 4061 895 4119 901
rect 4253 895 4311 901
rect 4445 895 4503 901
rect 2333 861 2345 895
rect 2525 861 2537 895
rect 2717 861 2729 895
rect 2909 861 2921 895
rect 3101 861 3113 895
rect 3293 861 3305 895
rect 3485 861 3497 895
rect 3677 861 3689 895
rect 3869 861 3881 895
rect 4061 861 4073 895
rect 4253 861 4265 895
rect 4445 861 4457 895
rect 2333 855 2391 861
rect 2525 855 2583 861
rect 2717 855 2775 861
rect 2909 855 2967 861
rect 3101 855 3159 861
rect 3293 855 3351 861
rect 3485 855 3543 861
rect 3677 855 3735 861
rect 3869 855 3927 861
rect 4061 855 4119 861
rect 4253 855 4311 861
rect 4445 855 4503 861
rect 2237 209 2295 215
rect 2429 209 2487 215
rect 2621 209 2679 215
rect 2813 209 2871 215
rect 3005 209 3063 215
rect 3197 209 3255 215
rect 3389 209 3447 215
rect 3581 209 3639 215
rect 3773 209 3831 215
rect 3965 209 4023 215
rect 4157 209 4215 215
rect 4349 209 4407 215
rect 2237 175 2249 209
rect 2429 175 2441 209
rect 2621 175 2633 209
rect 2813 175 2825 209
rect 3005 175 3017 209
rect 3197 175 3209 209
rect 3389 175 3401 209
rect 3581 175 3593 209
rect 3773 175 3785 209
rect 3965 175 3977 209
rect 4157 175 4169 209
rect 4349 175 4361 209
rect 2237 169 2295 175
rect 2429 169 2487 175
rect 2621 169 2679 175
rect 2813 169 2871 175
rect 3005 169 3063 175
rect 3197 169 3255 175
rect 3389 169 3447 175
rect 3581 169 3639 175
rect 3773 169 3831 175
rect 3965 169 4023 175
rect 4157 169 4215 175
rect 4349 169 4407 175
rect 2087 92 2102 126
rect 4638 73 4653 902
rect 4672 868 4707 902
rect 4672 73 4706 868
rect 4918 800 4976 806
rect 4918 766 4930 800
rect 4918 760 4976 766
rect 4822 156 4880 162
rect 5014 156 5072 162
rect 4822 122 4834 156
rect 5014 122 5026 156
rect 4822 116 4880 122
rect 5014 116 5072 122
rect 4672 39 4687 73
rect 5207 20 5222 902
rect 5241 20 5275 956
rect 5241 -14 5256 20
rect 5556 -33 5571 4206
rect 5590 4172 5625 4206
rect 5590 -33 5624 4172
rect 5886 1303 5920 1357
rect 5590 -67 5605 -33
rect 5905 -86 5920 1303
rect 5939 1269 5974 1303
rect 5939 -86 5973 1269
rect 6303 556 6337 610
rect 5939 -120 5954 -86
rect 6322 -139 6337 556
rect 6356 522 6391 556
rect 6356 -139 6390 522
rect 6602 454 6660 460
rect 6602 420 6614 454
rect 6602 414 6660 420
rect 6506 -56 6564 -50
rect 6698 -56 6756 -50
rect 6506 -90 6518 -56
rect 6698 -90 6710 -56
rect 6506 -96 6564 -90
rect 6698 -96 6756 -90
rect 6356 -173 6371 -139
use DAC  x1
timestamp 1752588718
transform 1 0 53 0 1 3436
box -2568 -3664 9162 4230
<< end >>
