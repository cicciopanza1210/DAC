magic
tech sky130A
magscale 1 2
timestamp 1753101330
<< error_p >>
rect 549 21896 550 22296
<< error_s >>
rect 7560 25589 7597 25590
rect 7885 25589 7914 25590
rect 7560 25380 7561 25589
rect 7913 25380 7914 25589
rect 8764 25359 8765 25626
rect 9231 25359 9232 25626
rect 10060 25621 10141 25622
rect 10429 25621 10462 25622
rect 10060 25385 10061 25621
rect 10461 25385 10462 25621
rect 11386 25391 11387 25628
rect 11787 25391 11788 25628
rect 11386 25390 11788 25391
rect 12840 25499 12911 25500
rect 13209 25499 13262 25500
rect 10060 25384 10462 25385
rect 8764 25358 9232 25359
rect 12840 25253 12841 25499
rect 13261 25253 13262 25499
rect 12840 25252 13262 25253
<< metal1 >>
rect 2284 26380 14727 26580
rect 234 21896 244 22296
rect 550 22184 560 22296
rect 2284 22184 2484 26380
rect 7526 25314 7536 25626
rect 7936 25314 7946 25626
rect 8744 25336 8754 25652
rect 9240 25336 9250 25652
rect 10022 25340 10032 25656
rect 10518 25340 10528 25656
rect 11342 25350 11352 25666
rect 11838 25350 11848 25666
rect 12808 25482 12818 25542
rect 7666 24888 7866 25314
rect 8914 24836 9114 25336
rect 10196 24748 10396 25340
rect 11494 24804 11694 25350
rect 11990 25282 12818 25482
rect 11990 24628 12190 25282
rect 12808 25226 12818 25282
rect 13304 25226 13314 25542
rect 14527 24467 14727 26380
rect 550 22108 3252 22184
rect 550 21896 560 22108
rect 3176 21970 3252 22108
rect 1012 20168 1022 20428
rect 1456 20376 1466 20428
rect 1642 20376 8548 20456
rect 1456 20252 8548 20376
rect 1456 20168 1466 20252
rect 1642 20228 8548 20252
<< via1 >>
rect 244 21896 550 22296
rect 7536 25314 7936 25626
rect 8754 25336 9240 25652
rect 10032 25340 10518 25656
rect 11352 25350 11838 25666
rect 12818 25226 13304 25542
rect 1022 20168 1456 20428
<< metal2 >>
rect 11352 25666 11456 25676
rect 11726 25666 11838 25676
rect 8754 25652 8826 25662
rect 9096 25652 9240 25662
rect 7536 25626 7624 25636
rect 7884 25626 7936 25636
rect 8754 25326 9240 25336
rect 10032 25656 10162 25666
rect 10432 25656 10518 25666
rect 11352 25340 11838 25350
rect 12818 25542 12916 25552
rect 13186 25542 13304 25552
rect 10032 25330 10518 25340
rect 7536 25304 7936 25314
rect 12818 25216 13304 25226
rect 244 22296 550 22306
rect 244 21886 550 21896
rect 890 20458 1144 20468
rect 1144 20428 1456 20438
rect 1144 20158 1456 20168
rect 890 20108 1144 20118
<< via2 >>
rect 7560 25380 7914 25590
rect 8764 25358 9232 25626
rect 10060 25384 10462 25622
rect 11386 25390 11788 25628
rect 12840 25252 13262 25500
rect 244 21896 550 22296
rect 890 20428 1144 20458
rect 890 20168 1022 20428
rect 1022 20168 1144 20428
rect 890 20118 1144 20168
<< metal3 >>
rect 8754 25626 9242 25631
rect 11376 25628 11798 25633
rect 7550 25590 7924 25595
rect 7550 25380 7560 25590
rect 7914 25380 7924 25590
rect 7550 25375 7924 25380
rect 8754 25358 8764 25626
rect 9232 25358 9242 25626
rect 10050 25622 10472 25627
rect 10050 25384 10060 25622
rect 10462 25384 10472 25622
rect 11376 25390 11386 25628
rect 11788 25390 11798 25628
rect 11376 25385 11798 25390
rect 12830 25500 13272 25505
rect 10050 25379 10472 25384
rect 8754 25353 9242 25358
rect 12830 25252 12840 25500
rect 13262 25252 13272 25500
rect 12830 25247 13272 25252
rect 234 22296 560 22301
rect 234 21896 244 22296
rect 550 21896 560 22296
rect 234 21891 560 21896
rect 880 20458 1154 20463
rect 880 20118 890 20458
rect 1144 20118 1154 20458
rect 880 20113 1154 20118
<< via3 >>
rect 7560 25380 7914 25590
rect 8764 25358 9232 25626
rect 10060 25384 10462 25622
rect 11386 25390 11788 25628
rect 12840 25252 13262 25500
rect 244 21896 550 22296
rect 890 20118 1144 20458
<< metal4 >>
rect 6134 44840 6194 45152
rect 6686 44840 6746 45152
rect 7238 44840 7298 45152
rect 7790 44840 7850 45152
rect 8342 44840 8402 45152
rect 8894 44840 8954 45152
rect 9446 44840 9506 45152
rect 9998 44840 10058 45152
rect 10550 44840 10610 45152
rect 11102 44840 11162 45152
rect 11654 44840 11714 45152
rect 12206 44840 12266 45152
rect 12758 44840 12818 45152
rect 13310 44840 13370 45152
rect 13862 44840 13922 45152
rect 14414 44840 14474 45152
rect 14966 44840 15026 45152
rect 15518 44840 15578 45152
rect 16070 44840 16130 45152
rect 16622 44840 16682 45152
rect 17174 44840 17234 45152
rect 17726 44840 17786 45152
rect 18278 44840 18338 45152
rect 18830 44840 18890 45152
rect 19382 44920 19442 45152
rect 19934 44920 19994 45152
rect 20486 44920 20546 45152
rect 21038 44920 21098 45152
rect 21590 44920 21650 45152
rect 22142 44920 22202 45152
rect 22694 44920 22754 45152
rect 23246 44920 23306 45152
rect 23798 44950 23858 45152
rect 24350 44950 24410 45152
rect 24902 44950 24962 45152
rect 25454 44950 25514 45152
rect 6134 44780 18926 44840
rect 6134 44152 6194 44780
rect 26006 44609 26066 45152
rect 7596 44319 26092 44609
rect 200 22296 600 44152
rect 800 43752 6256 44152
rect 200 21896 244 22296
rect 200 1000 600 21896
rect 800 20458 1200 43752
rect 7596 25590 7886 44319
rect 26558 44173 26618 45152
rect 8866 43891 26658 44173
rect 8866 27062 9148 43891
rect 27110 43353 27170 45152
rect 10140 43063 27173 43353
rect 8764 25626 9232 27062
rect 7560 25252 7914 25380
rect 10140 25622 10430 43063
rect 27662 42762 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 11428 42682 27775 42762
rect 11432 42472 27775 42682
rect 11432 27062 11722 42472
rect 12910 27598 30682 27898
rect 11386 25628 11788 27062
rect 12910 25500 13210 27598
rect 800 20118 890 20458
rect 1144 20118 1200 20458
rect 800 1000 1200 20118
rect 30382 8274 30682 27598
rect 30362 7920 30682 8274
rect 3314 0 3494 200
rect 7178 0 7358 200
rect 11042 0 11222 200
rect 14906 0 15086 200
rect 18770 0 18950 200
rect 22634 0 22814 200
rect 26498 0 26678 200
rect 30362 0 30542 7920
use DAC  DAC_0
timestamp 1752679897
transform 1 0 5578 0 1 22792
box -2462 -2574 9149 3152
<< labels >>
flabel metal4 200 1000 600 44152 1 FreeSans 1600 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 800 1000 1200 44152 1 FreeSans 1600 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
