magic
tech sky130A
magscale 1 2
timestamp 1751989567
<< error_p >>
rect -461 347 -403 353
rect -269 347 -211 353
rect -77 347 -19 353
rect 115 347 173 353
rect 307 347 365 353
rect 499 347 557 353
rect -461 313 -449 347
rect -269 313 -257 347
rect -77 313 -65 347
rect 115 313 127 347
rect 307 313 319 347
rect 499 313 511 347
rect -461 307 -403 313
rect -269 307 -211 313
rect -77 307 -19 313
rect 115 307 173 313
rect 307 307 365 313
rect 499 307 557 313
rect -557 -313 -499 -307
rect -365 -313 -307 -307
rect -173 -313 -115 -307
rect 19 -313 77 -307
rect 211 -313 269 -307
rect 403 -313 461 -307
rect -557 -347 -545 -313
rect -365 -347 -353 -313
rect -173 -347 -161 -313
rect 19 -347 31 -313
rect 211 -347 223 -313
rect 403 -347 415 -313
rect -557 -353 -499 -347
rect -365 -353 -307 -347
rect -173 -353 -115 -347
rect 19 -353 77 -347
rect 211 -353 269 -347
rect 403 -353 461 -347
<< pwell >>
rect -743 -485 743 485
<< nmoslvt >>
rect -546 -275 -510 275
rect -450 -275 -414 275
rect -354 -275 -318 275
rect -258 -275 -222 275
rect -162 -275 -126 275
rect -66 -275 -30 275
rect 30 -275 66 275
rect 126 -275 162 275
rect 222 -275 258 275
rect 318 -275 354 275
rect 414 -275 450 275
rect 510 -275 546 275
<< ndiff >>
rect -605 263 -546 275
rect -605 -263 -593 263
rect -559 -263 -546 263
rect -605 -275 -546 -263
rect -510 263 -450 275
rect -510 -263 -497 263
rect -463 -263 -450 263
rect -510 -275 -450 -263
rect -414 263 -354 275
rect -414 -263 -401 263
rect -367 -263 -354 263
rect -414 -275 -354 -263
rect -318 263 -258 275
rect -318 -263 -305 263
rect -271 -263 -258 263
rect -318 -275 -258 -263
rect -222 263 -162 275
rect -222 -263 -209 263
rect -175 -263 -162 263
rect -222 -275 -162 -263
rect -126 263 -66 275
rect -126 -263 -113 263
rect -79 -263 -66 263
rect -126 -275 -66 -263
rect -30 263 30 275
rect -30 -263 -17 263
rect 17 -263 30 263
rect -30 -275 30 -263
rect 66 263 126 275
rect 66 -263 79 263
rect 113 -263 126 263
rect 66 -275 126 -263
rect 162 263 222 275
rect 162 -263 175 263
rect 209 -263 222 263
rect 162 -275 222 -263
rect 258 263 318 275
rect 258 -263 271 263
rect 305 -263 318 263
rect 258 -275 318 -263
rect 354 263 414 275
rect 354 -263 367 263
rect 401 -263 414 263
rect 354 -275 414 -263
rect 450 263 510 275
rect 450 -263 463 263
rect 497 -263 510 263
rect 450 -275 510 -263
rect 546 263 605 275
rect 546 -263 559 263
rect 593 -263 605 263
rect 546 -275 605 -263
<< ndiffc >>
rect -593 -263 -559 263
rect -497 -263 -463 263
rect -401 -263 -367 263
rect -305 -263 -271 263
rect -209 -263 -175 263
rect -113 -263 -79 263
rect -17 -263 17 263
rect 79 -263 113 263
rect 175 -263 209 263
rect 271 -263 305 263
rect 367 -263 401 263
rect 463 -263 497 263
rect 559 -263 593 263
<< psubdiff >>
rect -707 415 -611 449
rect 611 415 707 449
rect -707 353 -673 415
rect 673 353 707 415
rect -707 -415 -673 -353
rect 673 -415 707 -353
rect -707 -449 -611 -415
rect 611 -449 707 -415
<< psubdiffcont >>
rect -611 415 611 449
rect -707 -353 -673 353
rect 673 -353 707 353
rect -611 -449 611 -415
<< poly >>
rect -465 347 -399 363
rect -465 313 -449 347
rect -415 313 -399 347
rect -546 275 -510 301
rect -465 297 -399 313
rect -273 347 -207 363
rect -273 313 -257 347
rect -223 313 -207 347
rect -450 275 -414 297
rect -354 275 -318 301
rect -273 297 -207 313
rect -81 347 -15 363
rect -81 313 -65 347
rect -31 313 -15 347
rect -258 275 -222 297
rect -162 275 -126 301
rect -81 297 -15 313
rect 111 347 177 363
rect 111 313 127 347
rect 161 313 177 347
rect -66 275 -30 297
rect 30 275 66 301
rect 111 297 177 313
rect 303 347 369 363
rect 303 313 319 347
rect 353 313 369 347
rect 126 275 162 297
rect 222 275 258 301
rect 303 297 369 313
rect 495 347 561 363
rect 495 313 511 347
rect 545 313 561 347
rect 318 275 354 297
rect 414 275 450 301
rect 495 297 561 313
rect 510 275 546 297
rect -546 -297 -510 -275
rect -561 -313 -495 -297
rect -450 -301 -414 -275
rect -354 -297 -318 -275
rect -561 -347 -545 -313
rect -511 -347 -495 -313
rect -561 -363 -495 -347
rect -369 -313 -303 -297
rect -258 -301 -222 -275
rect -162 -297 -126 -275
rect -369 -347 -353 -313
rect -319 -347 -303 -313
rect -369 -363 -303 -347
rect -177 -313 -111 -297
rect -66 -301 -30 -275
rect 30 -297 66 -275
rect -177 -347 -161 -313
rect -127 -347 -111 -313
rect -177 -363 -111 -347
rect 15 -313 81 -297
rect 126 -301 162 -275
rect 222 -297 258 -275
rect 15 -347 31 -313
rect 65 -347 81 -313
rect 15 -363 81 -347
rect 207 -313 273 -297
rect 318 -301 354 -275
rect 414 -297 450 -275
rect 207 -347 223 -313
rect 257 -347 273 -313
rect 207 -363 273 -347
rect 399 -313 465 -297
rect 510 -301 546 -275
rect 399 -347 415 -313
rect 449 -347 465 -313
rect 399 -363 465 -347
<< polycont >>
rect -449 313 -415 347
rect -257 313 -223 347
rect -65 313 -31 347
rect 127 313 161 347
rect 319 313 353 347
rect 511 313 545 347
rect -545 -347 -511 -313
rect -353 -347 -319 -313
rect -161 -347 -127 -313
rect 31 -347 65 -313
rect 223 -347 257 -313
rect 415 -347 449 -313
<< locali >>
rect -707 415 -611 449
rect 611 415 707 449
rect -707 353 -673 415
rect 673 353 707 415
rect -465 313 -449 347
rect -415 313 -399 347
rect -273 313 -257 347
rect -223 313 -207 347
rect -81 313 -65 347
rect -31 313 -15 347
rect 111 313 127 347
rect 161 313 177 347
rect 303 313 319 347
rect 353 313 369 347
rect 495 313 511 347
rect 545 313 561 347
rect -593 263 -559 279
rect -593 -279 -559 -263
rect -497 263 -463 279
rect -497 -279 -463 -263
rect -401 263 -367 279
rect -401 -279 -367 -263
rect -305 263 -271 279
rect -305 -279 -271 -263
rect -209 263 -175 279
rect -209 -279 -175 -263
rect -113 263 -79 279
rect -113 -279 -79 -263
rect -17 263 17 279
rect -17 -279 17 -263
rect 79 263 113 279
rect 79 -279 113 -263
rect 175 263 209 279
rect 175 -279 209 -263
rect 271 263 305 279
rect 271 -279 305 -263
rect 367 263 401 279
rect 367 -279 401 -263
rect 463 263 497 279
rect 463 -279 497 -263
rect 559 263 593 279
rect 559 -279 593 -263
rect -561 -347 -545 -313
rect -511 -347 -495 -313
rect -369 -347 -353 -313
rect -319 -347 -303 -313
rect -177 -347 -161 -313
rect -127 -347 -111 -313
rect 15 -347 31 -313
rect 65 -347 81 -313
rect 207 -347 223 -313
rect 257 -347 273 -313
rect 399 -347 415 -313
rect 449 -347 465 -313
rect -707 -415 -673 -353
rect 673 -415 707 -353
rect -707 -449 -611 -415
rect 611 -449 707 -415
<< viali >>
rect -449 313 -415 347
rect -257 313 -223 347
rect -65 313 -31 347
rect 127 313 161 347
rect 319 313 353 347
rect 511 313 545 347
rect -593 -263 -559 263
rect -497 -263 -463 263
rect -401 -263 -367 263
rect -305 -263 -271 263
rect -209 -263 -175 263
rect -113 -263 -79 263
rect -17 -263 17 263
rect 79 -263 113 263
rect 175 -263 209 263
rect 271 -263 305 263
rect 367 -263 401 263
rect 463 -263 497 263
rect 559 -263 593 263
rect -545 -347 -511 -313
rect -353 -347 -319 -313
rect -161 -347 -127 -313
rect 31 -347 65 -313
rect 223 -347 257 -313
rect 415 -347 449 -313
<< metal1 >>
rect -461 347 -403 353
rect -461 313 -449 347
rect -415 313 -403 347
rect -461 307 -403 313
rect -269 347 -211 353
rect -269 313 -257 347
rect -223 313 -211 347
rect -269 307 -211 313
rect -77 347 -19 353
rect -77 313 -65 347
rect -31 313 -19 347
rect -77 307 -19 313
rect 115 347 173 353
rect 115 313 127 347
rect 161 313 173 347
rect 115 307 173 313
rect 307 347 365 353
rect 307 313 319 347
rect 353 313 365 347
rect 307 307 365 313
rect 499 347 557 353
rect 499 313 511 347
rect 545 313 557 347
rect 499 307 557 313
rect -599 263 -553 275
rect -599 -263 -593 263
rect -559 -263 -553 263
rect -599 -275 -553 -263
rect -503 263 -457 275
rect -503 -263 -497 263
rect -463 -263 -457 263
rect -503 -275 -457 -263
rect -407 263 -361 275
rect -407 -263 -401 263
rect -367 -263 -361 263
rect -407 -275 -361 -263
rect -311 263 -265 275
rect -311 -263 -305 263
rect -271 -263 -265 263
rect -311 -275 -265 -263
rect -215 263 -169 275
rect -215 -263 -209 263
rect -175 -263 -169 263
rect -215 -275 -169 -263
rect -119 263 -73 275
rect -119 -263 -113 263
rect -79 -263 -73 263
rect -119 -275 -73 -263
rect -23 263 23 275
rect -23 -263 -17 263
rect 17 -263 23 263
rect -23 -275 23 -263
rect 73 263 119 275
rect 73 -263 79 263
rect 113 -263 119 263
rect 73 -275 119 -263
rect 169 263 215 275
rect 169 -263 175 263
rect 209 -263 215 263
rect 169 -275 215 -263
rect 265 263 311 275
rect 265 -263 271 263
rect 305 -263 311 263
rect 265 -275 311 -263
rect 361 263 407 275
rect 361 -263 367 263
rect 401 -263 407 263
rect 361 -275 407 -263
rect 457 263 503 275
rect 457 -263 463 263
rect 497 -263 503 263
rect 457 -275 503 -263
rect 553 263 599 275
rect 553 -263 559 263
rect 593 -263 599 263
rect 553 -275 599 -263
rect -557 -313 -499 -307
rect -557 -347 -545 -313
rect -511 -347 -499 -313
rect -557 -353 -499 -347
rect -365 -313 -307 -307
rect -365 -347 -353 -313
rect -319 -347 -307 -313
rect -365 -353 -307 -347
rect -173 -313 -115 -307
rect -173 -347 -161 -313
rect -127 -347 -115 -313
rect -173 -353 -115 -347
rect 19 -313 77 -307
rect 19 -347 31 -313
rect 65 -347 77 -313
rect 19 -353 77 -347
rect 211 -313 269 -307
rect 211 -347 223 -313
rect 257 -347 269 -313
rect 211 -353 269 -347
rect 403 -313 461 -307
rect 403 -347 415 -313
rect 449 -347 461 -313
rect 403 -353 461 -347
<< properties >>
string FIXED_BBOX -690 -432 690 432
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2.75 l 0.18 m 1 nf 12 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
