magic
tech sky130A
magscale 1 2
timestamp 1752767494
<< metal1 >>
rect 682 26926 692 27428
rect 1032 27268 1042 27428
rect 1032 27068 14541 27268
rect 1032 26926 1042 27068
rect 11076 26408 11086 26498
rect 11222 26473 11232 26498
rect 11222 26408 11237 26473
rect 7438 26196 7448 26318
rect 7710 26196 7720 26318
rect 7480 25636 7680 26196
rect 8642 26182 8652 26344
rect 8944 26182 8954 26344
rect 11107 26275 11237 26408
rect 8726 25556 8926 26182
rect 10000 26134 10010 26272
rect 10294 26134 10304 26272
rect 11107 26250 11238 26275
rect 11107 26248 11280 26250
rect 11107 26145 11506 26248
rect 10010 25484 10210 26134
rect 11306 25524 11506 26145
rect 11754 25940 11764 26126
rect 12082 25940 12092 26126
rect 11804 25348 12004 25940
rect 14341 25187 14541 27068
rect 2942 23232 2952 23246
rect 2930 23046 2952 23232
rect 3232 23046 3242 23246
rect 2930 22570 3130 23046
rect 7840 20938 8362 21166
rect 7840 20780 8068 20938
rect 7804 20562 7814 20780
rect 8076 20562 8086 20780
rect 18734 20564 18744 20806
rect 19208 20564 19218 20806
rect 18910 2914 19086 20564
rect 29466 8214 30078 8224
rect 29466 7214 30078 7224
rect 18910 2738 30324 2914
rect 30148 870 30324 2738
rect 30148 694 30530 870
rect 30354 586 30530 694
rect 30276 400 30286 586
rect 30654 400 30664 586
<< via1 >>
rect 692 26926 1032 27428
rect 11086 26408 11222 26498
rect 7448 26196 7710 26318
rect 8652 26182 8944 26344
rect 10010 26134 10294 26272
rect 11764 25940 12082 26126
rect 2952 23046 3232 23246
rect 7814 20562 8076 20780
rect 18744 20564 19208 20806
rect 29466 7224 30078 8214
rect 30286 400 30654 586
<< metal2 >>
rect 692 27428 1032 27438
rect 692 26916 1032 26926
rect 11086 26498 11222 26508
rect 11086 26398 11222 26408
rect 8652 26344 8944 26354
rect 7448 26318 7710 26328
rect 7448 26186 7710 26196
rect 8652 26172 8944 26182
rect 10010 26272 10294 26282
rect 10010 26124 10294 26134
rect 11764 26126 12082 26136
rect 12082 25976 19033 26082
rect 11764 25930 12082 25940
rect 1374 23564 1910 23574
rect 1910 23173 1935 23357
rect 2952 23246 3232 23256
rect 1910 23118 2952 23173
rect 1910 22920 1935 23118
rect 2952 23036 3232 23046
rect 1374 22910 1935 22920
rect 1873 22884 1935 22910
rect 18927 20816 19033 25976
rect 18744 20806 19208 20816
rect 7814 20780 8076 20790
rect 7814 20552 8076 20562
rect 18744 20554 19208 20564
rect 7832 20287 8076 20552
rect 7832 20152 28748 20287
rect 7885 20148 28748 20152
rect 28609 7759 28748 20148
rect 29456 8212 29466 8214
rect 29448 7759 29466 8212
rect 28609 7625 29466 7759
rect 28609 7623 28748 7625
rect 29448 7234 29466 7625
rect 29456 7224 29466 7234
rect 30078 7224 30088 8214
rect 30286 586 30654 596
rect 30286 390 30654 400
<< via2 >>
rect 692 26926 1032 27428
rect 11086 26408 11222 26498
rect 7448 26196 7710 26318
rect 8652 26182 8944 26344
rect 10010 26134 10294 26272
rect 1374 22920 1910 23564
rect 29466 7224 30078 8214
rect 30286 400 30654 586
<< metal3 >>
rect 25314 43234 25324 43594
rect 25728 43527 25738 43594
rect 27956 43527 27966 43744
rect 25728 43310 27966 43527
rect 25728 43234 25738 43310
rect 27956 43210 27966 43310
rect 28490 43210 28500 43744
rect 682 27428 1042 27433
rect 682 26926 692 27428
rect 1032 26926 1042 27428
rect 682 26921 1042 26926
rect 11076 26498 11232 26503
rect 11076 26408 11086 26498
rect 11222 26408 11232 26498
rect 11076 26403 11232 26408
rect 8642 26344 8954 26349
rect 7438 26318 7720 26323
rect 7438 26196 7448 26318
rect 7710 26196 7720 26318
rect 7438 26191 7720 26196
rect 8642 26182 8652 26344
rect 8944 26182 8954 26344
rect 8642 26177 8954 26182
rect 10000 26272 10304 26277
rect 10000 26134 10010 26272
rect 10294 26134 10304 26272
rect 10000 26129 10304 26134
rect 1364 23564 1920 23569
rect 1364 23558 1374 23564
rect 1162 22914 1172 23558
rect 1910 22920 1920 23564
rect 1708 22915 1920 22920
rect 1708 22914 1718 22915
rect 29461 8214 30083 8224
rect 29461 7224 29466 8214
rect 30078 7224 30083 8214
rect 29461 7214 30083 7224
rect 30276 586 30664 591
rect 30276 400 30286 586
rect 30654 400 30664 586
rect 30276 395 30664 400
<< via3 >>
rect 25324 43234 25728 43594
rect 27966 43210 28490 43744
rect 692 26926 1032 27428
rect 11086 26408 11222 26498
rect 7448 26196 7710 26318
rect 8652 26182 8944 26344
rect 10010 26134 10294 26272
rect 1172 22920 1374 23558
rect 1374 22920 1708 23558
rect 1172 22914 1708 22920
rect 29466 7224 30078 8214
rect 30286 400 30654 586
<< metal4 >>
rect 200 27380 600 44152
rect 6134 43543 6194 45152
rect 6686 43543 6746 45152
rect 7238 43543 7298 45152
rect 7790 43543 7850 45152
rect 8342 43543 8402 45152
rect 8894 43543 8954 45152
rect 9446 43543 9506 45152
rect 9998 43543 10058 45152
rect 10550 43543 10610 45152
rect 11102 43543 11162 45152
rect 11654 43543 11714 45152
rect 12206 43543 12266 45152
rect 12758 43543 12818 45152
rect 13310 43543 13370 45152
rect 13862 43543 13922 45152
rect 14414 43543 14474 45152
rect 14966 43543 15026 45152
rect 15518 43543 15578 45152
rect 16070 43543 16130 45152
rect 16622 43543 16682 45152
rect 17174 43543 17234 45152
rect 17726 43543 17786 45152
rect 18278 43543 18338 45152
rect 18830 43543 18890 45152
rect 19382 43543 19442 45152
rect 19934 43543 19994 45152
rect 20486 43543 20546 45152
rect 21038 43543 21098 45152
rect 21590 43543 21650 45152
rect 22142 43543 22202 45152
rect 22694 43543 22754 45152
rect 23246 43543 23306 45152
rect 23798 43543 23858 45152
rect 24350 43543 24410 45152
rect 24902 43543 24962 45152
rect 25454 43774 25514 45152
rect 25096 43714 25514 43774
rect 25096 43543 25156 43714
rect 25323 43594 25729 43595
rect 25323 43543 25324 43594
rect 6104 43326 25324 43543
rect 25323 43234 25324 43326
rect 25728 43234 25729 43594
rect 25323 43233 25729 43234
rect 26006 42238 26066 45152
rect 7738 42178 26066 42238
rect 691 27428 1033 27429
rect 691 27380 692 27428
rect 200 26980 692 27380
rect 200 23438 600 26980
rect 691 26926 692 26980
rect 1032 26926 1033 27428
rect 691 26925 1033 26926
rect 7738 26456 7798 42178
rect 26558 41902 26618 45152
rect 9290 41842 26618 41902
rect 9296 26708 9356 41842
rect 27110 41574 27170 45152
rect 7564 26396 7798 26456
rect 7564 26319 7624 26396
rect 7738 26390 7798 26396
rect 8790 26648 9356 26708
rect 8790 26345 8850 26648
rect 9296 26638 9356 26648
rect 10316 41514 27170 41574
rect 10316 26644 10376 41514
rect 27662 41288 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 27965 43744 28491 43745
rect 27965 43210 27966 43744
rect 28490 43694 28491 43744
rect 28490 43294 32014 43694
rect 28490 43210 28491 43294
rect 27965 43209 28491 43210
rect 10084 26600 10376 26644
rect 11126 41228 27722 41288
rect 10084 26540 10378 26600
rect 8651 26344 8945 26345
rect 7447 26318 7711 26319
rect 7447 26196 7448 26318
rect 7710 26196 7711 26318
rect 7447 26195 7711 26196
rect 8651 26182 8652 26344
rect 8944 26182 8945 26344
rect 10084 26273 10220 26540
rect 11126 26499 11186 41228
rect 11085 26498 11223 26499
rect 11085 26408 11086 26498
rect 11222 26408 11223 26498
rect 11085 26407 11223 26408
rect 8651 26181 8945 26182
rect 10009 26272 10295 26273
rect 10009 26134 10010 26272
rect 10294 26134 10295 26272
rect 10009 26133 10295 26134
rect 1171 23558 1709 23559
rect 1171 23438 1172 23558
rect 200 23038 1172 23438
rect 200 1000 600 23038
rect 1171 22914 1172 23038
rect 1708 22914 1709 23558
rect 1171 22913 1709 22914
rect 29465 8214 30079 8215
rect 29465 7224 29466 8214
rect 30078 7954 30079 8214
rect 31614 7954 32014 43294
rect 30078 7554 32014 7954
rect 30078 7224 30079 7554
rect 29465 7223 30079 7224
rect 30285 586 30655 587
rect 30285 400 30286 586
rect 30654 400 30655 586
rect 31614 542 32014 7554
rect 30285 399 30655 400
rect 3314 0 3494 212
rect 7178 0 7358 212
rect 11042 0 11222 212
rect 14906 0 15086 206
rect 18770 0 18950 206
rect 22634 0 22814 206
rect 26498 0 26678 206
rect 30362 0 30542 399
use untitled-3  untitled-3_0
timestamp 1752761699
transform 1 0 5339 0 1 20076
box -2409 862 9202 6588
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 11042 0 11222 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 7178 0 7358 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 3314 0 3494 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 1600 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 31614 542 32014 43694 1 FreeSans 1600 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
