* SPICE3 file created from tt_um_DAC1.ext - technology: sky130A

X0 VGND DAC_0/m1_n1165_n912# DAC_0/m1_n1165_n912# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.78765 pd=5.93 as=0.4005 ps=2.97 w=2.67 l=0.18
X1 VGND DAC_0/m1_n1165_n912# DAC_0/m1_n1165_n912# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.4005 pd=2.97 as=0.78765 ps=5.93 w=2.67 l=0.18
X2 DAC_0/m1_n1165_n912# DAC_0/m1_n1165_n912# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.4005 pd=2.97 as=0.4005 ps=2.97 w=2.67 l=0.18
X3 VGND DAC_0/m1_n1165_n912# DAC_0/m1_1348_n950# VGND sky130_fd_pr__nfet_01v8_lvt ad=20.8983 pd=154.48 as=2.77865 ps=21.06 w=2.67 l=0.18
X4 VGND DAC_0/m1_n1165_n912# DAC_0/m1_1348_n950# VGND sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2.67 l=0.18
X5 DAC_0/m1_1348_n950# DAC_0/m1_n1165_n912# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2.67 l=0.18
X6 DAC_0/m1_2538_n916# DAC_0/m1_n1165_n912# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.4005 pd=2.97 as=0.4005 ps=2.97 w=2.67 l=0.18
X7 VGND DAC_0/m1_n1165_n912# DAC_0/m1_2538_n916# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.4005 pd=2.97 as=0.78765 ps=5.93 w=2.67 l=0.18
X8 DAC_0/m1_2538_n916# DAC_0/m1_n1165_n912# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.78765 pd=5.93 as=0.4005 ps=2.97 w=2.67 l=0.18
X9 DAC_0/m1_2538_n916# DAC_0/m1_n1165_n912# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.4005 pd=2.97 as=0.4005 ps=2.97 w=2.67 l=0.18
X10 VGND DAC_0/m1_n1165_n912# DAC_0/m1_2538_n916# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.4005 pd=2.97 as=0.4005 ps=2.97 w=2.67 l=0.18
X11 VGND DAC_0/m1_n1165_n912# DAC_0/m1_2538_n916# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.4005 pd=2.97 as=0.4005 ps=2.97 w=2.67 l=0.18
X12 DAC_0/m1_n1797_2673# VDPWR VGND sky130_fd_pr__res_xhigh_po_0p35 l=16
X13 ua[0] VDPWR VGND sky130_fd_pr__res_xhigh_po_0p69 l=1.75
X14 DAC_0/m1_5188_872# DAC_0/m1_n1165_n912# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X15 VGND DAC_0/m1_n1165_n912# DAC_0/m1_5188_872# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X16 VGND DAC_0/m1_n1165_n912# DAC_0/m1_5188_872# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X17 DAC_0/m1_5188_872# DAC_0/m1_n1165_n912# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X18 DAC_0/m1_5188_872# DAC_0/m1_n1165_n912# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X19 VGND DAC_0/m1_n1165_n912# DAC_0/m1_5188_872# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X20 VGND DAC_0/m1_n1165_n912# DAC_0/m1_5188_872# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.8496 ps=6.35 w=2.88 l=0.18
X21 DAC_0/m1_5188_872# DAC_0/m1_n1165_n912# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X22 DAC_0/m1_5188_872# DAC_0/m1_n1165_n912# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X23 VGND DAC_0/m1_n1165_n912# DAC_0/m1_5188_872# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X24 VGND DAC_0/m1_n1165_n912# DAC_0/m1_5188_872# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X25 VGND DAC_0/m1_n1165_n912# DAC_0/m1_5188_872# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X26 DAC_0/m1_5188_872# DAC_0/m1_n1165_n912# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.8496 pd=6.35 as=0.432 ps=3.18 w=2.88 l=0.18
X27 DAC_0/m1_5188_872# DAC_0/m1_n1165_n912# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X28 DAC_0/m1_5188_872# DAC_0/m1_n1165_n912# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X29 DAC_0/m1_5188_872# DAC_0/m1_n1165_n912# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X30 VGND DAC_0/m1_n1165_n912# DAC_0/m1_5188_872# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X31 VGND DAC_0/m1_n1165_n912# DAC_0/m1_5188_872# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X32 DAC_0/m1_5188_872# DAC_0/m1_n1165_n912# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X33 VGND DAC_0/m1_n1165_n912# DAC_0/m1_5188_872# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X34 VGND DAC_0/m1_n1165_n912# DAC_0/m1_5188_872# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X35 DAC_0/m1_5188_872# DAC_0/m1_n1165_n912# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X36 DAC_0/m1_5188_872# DAC_0/m1_n1165_n912# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X37 VGND DAC_0/m1_n1165_n912# DAC_0/m1_5188_872# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.432 pd=3.18 as=0.432 ps=3.18 w=2.88 l=0.18
X38 VGND DAC_0/m1_n1165_n912# DAC_0/m1_3770_n1012# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.4125 pd=3.05 as=0.4125 ps=3.05 w=2.75 l=0.18
X39 VGND DAC_0/m1_n1165_n912# DAC_0/m1_3770_n1012# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.4125 pd=3.05 as=0.4125 ps=3.05 w=2.75 l=0.18
X40 DAC_0/m1_3770_n1012# DAC_0/m1_n1165_n912# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.4125 pd=3.05 as=0.4125 ps=3.05 w=2.75 l=0.18
X41 DAC_0/m1_3770_n1012# DAC_0/m1_n1165_n912# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.4125 pd=3.05 as=0.4125 ps=3.05 w=2.75 l=0.18
X42 VGND DAC_0/m1_n1165_n912# DAC_0/m1_3770_n1012# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.4125 pd=3.05 as=0.81125 ps=6.09 w=2.75 l=0.18
X43 VGND DAC_0/m1_n1165_n912# DAC_0/m1_3770_n1012# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.4125 pd=3.05 as=0.4125 ps=3.05 w=2.75 l=0.18
X44 DAC_0/m1_3770_n1012# DAC_0/m1_n1165_n912# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.4125 pd=3.05 as=0.4125 ps=3.05 w=2.75 l=0.18
X45 DAC_0/m1_3770_n1012# DAC_0/m1_n1165_n912# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.81125 pd=6.09 as=0.4125 ps=3.05 w=2.75 l=0.18
X46 VGND DAC_0/m1_n1165_n912# DAC_0/m1_3770_n1012# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.4125 pd=3.05 as=0.4125 ps=3.05 w=2.75 l=0.18
X47 DAC_0/m1_3770_n1012# DAC_0/m1_n1165_n912# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.4125 pd=3.05 as=0.4125 ps=3.05 w=2.75 l=0.18
X48 DAC_0/m1_3770_n1012# DAC_0/m1_n1165_n912# VGND VGND sky130_fd_pr__nfet_01v8_lvt ad=0.4125 pd=3.05 as=0.4125 ps=3.05 w=2.75 l=0.18
X49 VGND DAC_0/m1_n1165_n912# DAC_0/m1_3770_n1012# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.4125 pd=3.05 as=0.4125 ps=3.05 w=2.75 l=0.18
X50 DAC_0/m1_1348_n950# ui_in[3] ua[0] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.59 pd=4.59 as=0.3 ps=2.3 w=2 l=0.18
X51 DAC_0/m1_1348_n950# ui_in[3] ua[0] VGND sky130_fd_pr__nfet_01v8_lvt ad=0.3 pd=2.3 as=0.59 ps=4.59 w=2 l=0.18
X52 ua[0] ui_in[3] DAC_0/m1_1348_n950# VGND sky130_fd_pr__nfet_01v8_lvt ad=0.3 pd=2.3 as=0.3 ps=2.3 w=2 l=0.18
X53 DAC_0/m1_n1797_2673# DAC_0/m1_n1165_n912# VGND sky130_fd_pr__res_xhigh_po_0p35 l=16
X54 DAC_0/m1_2538_n916# ui_in[2] ua[0] VGND sky130_fd_pr__nfet_01v8_lvt ad=4.3673 pd=32.93 as=4.76 ps=36.76 w=2 l=0.18
X55 DAC_0/m1_2538_n916# ui_in[2] ua[0] VGND sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2 l=0.18
X56 ua[0] ui_in[2] DAC_0/m1_2538_n916# VGND sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2 l=0.18
X57 DAC_0/m1_3770_n1012# ui_in[1] ua[0] VGND sky130_fd_pr__nfet_01v8_lvt ad=6.9375 pd=51.87 as=0 ps=0 w=2 l=0.18
X58 DAC_0/m1_3770_n1012# ui_in[1] ua[0] VGND sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2 l=0.18
X59 ua[0] ui_in[1] DAC_0/m1_3770_n1012# VGND sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2 l=0.18
X60 DAC_0/m1_5188_872# ui_in[0] ua[0] VGND sky130_fd_pr__nfet_01v8_lvt ad=12.3932 pd=91.85 as=0 ps=0 w=2 l=0.18
X61 DAC_0/m1_5188_872# ui_in[0] ua[0] VGND sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2 l=0.18
X62 ua[0] ui_in[0] DAC_0/m1_5188_872# VGND sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=2 l=0.18
C0 ui_in[0] ui_in[1] 5.457032f
C1 ui_in[1] ui_in[2] 4.223191f
C2 ui_in[2] ui_in[3] 8.091054f
C3 DAC_0/m1_5188_872# DAC_0/m1_n1165_n912# 2.419775f
C4 ui_in[0] VGND 12.856084f
C5 ui_in[1] VGND 8.950926f
C6 ui_in[2] VGND 9.215423f
C7 ua[0] VGND 25.7654f
C8 ui_in[3] VGND 15.420452f
C9 DAC_0/m1_3770_n1012# VGND 7.532216f **FLOATING
C10 DAC_0/m1_5188_872# VGND 13.893605f **FLOATING
C11 VDPWR VGND 31.084164f
C12 DAC_0/m1_2538_n916# VGND 4.484244f **FLOATING
C13 DAC_0/m1_1348_n950# VGND 2.994625f **FLOATING
C14 DAC_0/m1_n1165_n912# VGND 23.264309f **FLOATING
