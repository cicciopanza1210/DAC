magic
tech sky130A
magscale 1 2
timestamp 1751989567
<< error_p >>
rect -173 339 -115 345
rect 19 339 77 345
rect 211 339 269 345
rect -173 305 -161 339
rect 19 305 31 339
rect 211 305 223 339
rect -173 299 -115 305
rect 19 299 77 305
rect 211 299 269 305
rect -269 -305 -211 -299
rect -77 -305 -19 -299
rect 115 -305 173 -299
rect -269 -339 -257 -305
rect -77 -339 -65 -305
rect 115 -339 127 -305
rect -269 -345 -211 -339
rect -77 -345 -19 -339
rect 115 -345 173 -339
<< pwell >>
rect -455 -477 455 477
<< nmoslvt >>
rect -258 -267 -222 267
rect -162 -267 -126 267
rect -66 -267 -30 267
rect 30 -267 66 267
rect 126 -267 162 267
rect 222 -267 258 267
<< ndiff >>
rect -317 255 -258 267
rect -317 -255 -305 255
rect -271 -255 -258 255
rect -317 -267 -258 -255
rect -222 255 -162 267
rect -222 -255 -209 255
rect -175 -255 -162 255
rect -222 -267 -162 -255
rect -126 255 -66 267
rect -126 -255 -113 255
rect -79 -255 -66 255
rect -126 -267 -66 -255
rect -30 255 30 267
rect -30 -255 -17 255
rect 17 -255 30 255
rect -30 -267 30 -255
rect 66 255 126 267
rect 66 -255 79 255
rect 113 -255 126 255
rect 66 -267 126 -255
rect 162 255 222 267
rect 162 -255 175 255
rect 209 -255 222 255
rect 162 -267 222 -255
rect 258 255 317 267
rect 258 -255 271 255
rect 305 -255 317 255
rect 258 -267 317 -255
<< ndiffc >>
rect -305 -255 -271 255
rect -209 -255 -175 255
rect -113 -255 -79 255
rect -17 -255 17 255
rect 79 -255 113 255
rect 175 -255 209 255
rect 271 -255 305 255
<< psubdiff >>
rect -419 407 -323 441
rect 323 407 419 441
rect -419 345 -385 407
rect 385 345 419 407
rect -419 -407 -385 -345
rect 385 -407 419 -345
rect -419 -441 -323 -407
rect 323 -441 419 -407
<< psubdiffcont >>
rect -323 407 323 441
rect -419 -345 -385 345
rect 385 -345 419 345
rect -323 -441 323 -407
<< poly >>
rect -177 339 -111 355
rect -177 305 -161 339
rect -127 305 -111 339
rect -258 267 -222 293
rect -177 289 -111 305
rect 15 339 81 355
rect 15 305 31 339
rect 65 305 81 339
rect -162 267 -126 289
rect -66 267 -30 293
rect 15 289 81 305
rect 207 339 273 355
rect 207 305 223 339
rect 257 305 273 339
rect 30 267 66 289
rect 126 267 162 293
rect 207 289 273 305
rect 222 267 258 289
rect -258 -289 -222 -267
rect -273 -305 -207 -289
rect -162 -293 -126 -267
rect -66 -289 -30 -267
rect -273 -339 -257 -305
rect -223 -339 -207 -305
rect -273 -355 -207 -339
rect -81 -305 -15 -289
rect 30 -293 66 -267
rect 126 -289 162 -267
rect -81 -339 -65 -305
rect -31 -339 -15 -305
rect -81 -355 -15 -339
rect 111 -305 177 -289
rect 222 -293 258 -267
rect 111 -339 127 -305
rect 161 -339 177 -305
rect 111 -355 177 -339
<< polycont >>
rect -161 305 -127 339
rect 31 305 65 339
rect 223 305 257 339
rect -257 -339 -223 -305
rect -65 -339 -31 -305
rect 127 -339 161 -305
<< locali >>
rect -419 407 -323 441
rect 323 407 419 441
rect -419 345 -385 407
rect 385 345 419 407
rect -177 305 -161 339
rect -127 305 -111 339
rect 15 305 31 339
rect 65 305 81 339
rect 207 305 223 339
rect 257 305 273 339
rect -305 255 -271 271
rect -305 -271 -271 -255
rect -209 255 -175 271
rect -209 -271 -175 -255
rect -113 255 -79 271
rect -113 -271 -79 -255
rect -17 255 17 271
rect -17 -271 17 -255
rect 79 255 113 271
rect 79 -271 113 -255
rect 175 255 209 271
rect 175 -271 209 -255
rect 271 255 305 271
rect 271 -271 305 -255
rect -273 -339 -257 -305
rect -223 -339 -207 -305
rect -81 -339 -65 -305
rect -31 -339 -15 -305
rect 111 -339 127 -305
rect 161 -339 177 -305
rect -419 -407 -385 -345
rect 385 -407 419 -345
rect -419 -441 -323 -407
rect 323 -441 419 -407
<< viali >>
rect -161 305 -127 339
rect 31 305 65 339
rect 223 305 257 339
rect -305 -255 -271 255
rect -209 -255 -175 255
rect -113 -255 -79 255
rect -17 -255 17 255
rect 79 -255 113 255
rect 175 -255 209 255
rect 271 -255 305 255
rect -257 -339 -223 -305
rect -65 -339 -31 -305
rect 127 -339 161 -305
<< metal1 >>
rect -173 339 -115 345
rect -173 305 -161 339
rect -127 305 -115 339
rect -173 299 -115 305
rect 19 339 77 345
rect 19 305 31 339
rect 65 305 77 339
rect 19 299 77 305
rect 211 339 269 345
rect 211 305 223 339
rect 257 305 269 339
rect 211 299 269 305
rect -311 255 -265 267
rect -311 -255 -305 255
rect -271 -255 -265 255
rect -311 -267 -265 -255
rect -215 255 -169 267
rect -215 -255 -209 255
rect -175 -255 -169 255
rect -215 -267 -169 -255
rect -119 255 -73 267
rect -119 -255 -113 255
rect -79 -255 -73 255
rect -119 -267 -73 -255
rect -23 255 23 267
rect -23 -255 -17 255
rect 17 -255 23 255
rect -23 -267 23 -255
rect 73 255 119 267
rect 73 -255 79 255
rect 113 -255 119 255
rect 73 -267 119 -255
rect 169 255 215 267
rect 169 -255 175 255
rect 209 -255 215 255
rect 169 -267 215 -255
rect 265 255 311 267
rect 265 -255 271 255
rect 305 -255 311 255
rect 265 -267 311 -255
rect -269 -305 -211 -299
rect -269 -339 -257 -305
rect -223 -339 -211 -305
rect -269 -345 -211 -339
rect -77 -305 -19 -299
rect -77 -339 -65 -305
rect -31 -339 -19 -305
rect -77 -345 -19 -339
rect 115 -305 173 -299
rect 115 -339 127 -305
rect 161 -339 173 -305
rect 115 -345 173 -339
<< properties >>
string FIXED_BBOX -402 -424 402 424
string gencell sky130_fd_pr__nfet_01v8_lvt
string library sky130
string parameters w 2.6666666666666665 l 0.18 m 1 nf 6 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
