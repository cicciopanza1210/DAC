magic
tech sky130A
magscale 1 2
timestamp 1752679897
<< viali >>
rect 6890 1554 8168 1618
rect 5478 696 5860 742
rect 1632 630 2008 680
rect 2832 650 3214 696
rect 4164 644 4546 690
rect -1824 -1190 -1656 -1132
rect -1232 -1192 -1064 -1134
rect 138 -1580 516 -1522
rect 1616 -1602 1990 -1550
rect 2742 -1568 3414 -1516
rect 3978 -1686 5220 -1634
rect 5760 -1720 8160 -1666
<< metal1 >>
rect -1797 2673 -1003 2867
rect 2088 2124 2302 2324
rect 2088 2048 2288 2124
rect 2082 1916 2092 2048
rect 2288 1916 2298 2048
rect 3334 2044 3536 2244
rect 3334 1936 3534 2044
rect 4618 1936 4818 2172
rect 5914 2012 6116 2212
rect 5914 1972 6114 2012
rect 3334 1906 3378 1936
rect 3338 1856 3378 1906
rect 3498 1856 3538 1936
rect 4614 1916 4818 1936
rect 4614 1904 4676 1916
rect 3338 1846 3538 1856
rect 4616 1836 4676 1904
rect 4796 1858 4818 1916
rect 5912 1946 6114 1972
rect 5912 1866 5958 1946
rect 6078 1896 6114 1946
rect 6078 1866 6112 1896
rect 4796 1836 4816 1858
rect 5912 1848 6112 1866
rect 6412 1836 6612 2036
rect 8949 1840 9149 1875
rect 4616 1820 4816 1836
rect 6471 1762 6554 1836
rect 1416 1718 7188 1762
rect 1416 1134 1460 1718
rect 2058 1546 2068 1674
rect 2294 1546 2304 1674
rect 2154 1320 2218 1546
rect 1708 1256 2218 1320
rect 1638 1134 1648 1144
rect 1408 1090 1648 1134
rect 1638 1084 1648 1090
rect 1700 1084 1710 1144
rect 1653 1048 1708 1084
rect 1836 1082 1846 1142
rect 1898 1082 1908 1142
rect 1390 892 1400 902
rect 982 -356 992 -302
rect 671 -407 992 -356
rect 671 -439 722 -407
rect -127 -489 723 -439
rect 982 -488 992 -407
rect 1152 -488 1162 -302
rect -2462 -942 -1682 -742
rect -127 -870 -77 -489
rect 671 -491 723 -489
rect 673 -786 723 -491
rect 132 -814 726 -786
rect 144 -870 154 -868
rect -1165 -912 154 -870
rect -150 -920 154 -912
rect 144 -922 154 -920
rect 214 -922 224 -868
rect 338 -916 348 -862
rect 408 -916 418 -862
rect -1836 -1132 -1644 -1126
rect -1836 -1190 -1824 -1132
rect -1656 -1190 -1644 -1132
rect -1836 -1196 -1644 -1190
rect -1244 -1134 -1052 -1128
rect -1244 -1192 -1232 -1134
rect -1064 -1192 -1052 -1134
rect -1244 -1194 -1052 -1192
rect -1824 -1224 -1656 -1196
rect -1280 -1198 -1052 -1194
rect -1280 -1224 -1068 -1198
rect -1824 -1232 -1068 -1224
rect -1802 -1268 -1068 -1232
rect -1802 -1289 -70 -1268
rect -1802 -1304 -35 -1289
rect -1802 -1334 -104 -1304
rect -1110 -1374 -104 -1334
rect -40 -1374 -30 -1304
rect 240 -1366 250 -1312
rect 310 -1366 320 -1312
rect 434 -1362 444 -1308
rect 504 -1362 514 -1308
rect -1110 -1500 -50 -1374
rect 698 -1432 726 -814
rect 782 -878 792 -780
rect 898 -878 908 -780
rect 158 -1460 726 -1432
rect -106 -1820 -50 -1500
rect 126 -1522 528 -1516
rect 126 -1580 138 -1522
rect 516 -1580 528 -1522
rect 126 -1586 528 -1580
rect 158 -1820 478 -1586
rect 816 -1820 872 -878
rect 1348 -898 1400 892
rect 1466 832 1476 902
rect 1740 828 1750 888
rect 1802 828 1812 888
rect 1932 834 1942 894
rect 1994 834 2004 894
rect 2154 790 2218 1256
rect 2625 1176 2667 1718
rect 3408 1660 3468 1674
rect 3366 1554 3376 1660
rect 3504 1554 3514 1660
rect 3408 1322 3468 1554
rect 2834 1262 3490 1322
rect 2834 1176 2844 1182
rect 2620 1134 2844 1176
rect 2834 1128 2844 1134
rect 2904 1128 2914 1182
rect 3032 1132 3042 1186
rect 3102 1132 3112 1186
rect 2546 906 2556 908
rect 1598 726 2218 790
rect 2539 848 2556 906
rect 2630 848 2640 908
rect 2936 852 2946 906
rect 3006 852 3016 906
rect 3128 850 3138 904
rect 3198 850 3208 904
rect 1620 680 2020 686
rect 1620 630 1632 680
rect 2008 630 2020 680
rect 1620 624 2020 630
rect 1630 584 2012 624
rect 1648 486 2008 584
rect 1648 480 1774 486
rect 1764 410 1774 480
rect 1850 480 2008 486
rect 1850 410 1860 480
rect 2168 -424 2178 -358
rect 2250 -424 2260 -358
rect 2195 -802 2237 -424
rect 1624 -844 2250 -802
rect 1348 -904 1490 -898
rect 1620 -904 1630 -902
rect 1348 -950 1630 -904
rect 1416 -954 1630 -950
rect 1620 -956 1630 -954
rect 1690 -956 1700 -902
rect 1814 -954 1824 -900
rect 1884 -954 1894 -900
rect 1342 -1422 1352 -1332
rect 1442 -1422 1452 -1332
rect 1716 -1396 1726 -1342
rect 1786 -1396 1796 -1342
rect 1910 -1394 1920 -1340
rect 1980 -1394 1990 -1340
rect 1368 -1820 1424 -1422
rect 2195 -1461 2237 -844
rect 2539 -866 2588 848
rect 3408 790 3468 1262
rect 3948 1198 3990 1718
rect 4668 1586 4678 1674
rect 4802 1586 4812 1674
rect 4722 1308 4770 1586
rect 4178 1260 4770 1308
rect 4170 1198 4180 1206
rect 3948 1156 4180 1198
rect 4170 1152 4180 1156
rect 4240 1152 4250 1206
rect 4364 1154 4374 1208
rect 4434 1154 4444 1208
rect 3896 883 3906 900
rect 2866 730 3468 790
rect 3773 833 3906 883
rect 2820 696 3226 702
rect 2820 650 2832 696
rect 3214 650 3226 696
rect 2820 644 3226 650
rect 2832 606 3214 644
rect 2848 474 3208 606
rect 2980 398 2990 474
rect 3066 398 3076 474
rect 3530 -426 3540 -360
rect 3612 -426 3622 -360
rect 3559 -772 3589 -426
rect 2756 -802 3590 -772
rect 2742 -866 2752 -864
rect 2538 -916 2752 -866
rect 2742 -918 2752 -916
rect 2812 -918 2822 -864
rect 2938 -916 2948 -862
rect 3008 -916 3018 -862
rect 3130 -912 3140 -858
rect 3200 -912 3210 -858
rect 3322 -912 3332 -858
rect 3392 -912 3402 -858
rect 2452 -1384 2462 -1294
rect 2552 -1384 2562 -1294
rect 2842 -1362 2852 -1308
rect 2912 -1362 2922 -1308
rect 3034 -1360 3044 -1306
rect 3104 -1360 3114 -1306
rect 3228 -1354 3238 -1300
rect 3298 -1354 3308 -1300
rect 1589 -1503 2237 -1461
rect 1604 -1550 2002 -1544
rect 1604 -1602 1616 -1550
rect 1990 -1602 2002 -1550
rect 1604 -1608 2002 -1602
rect 1652 -1820 1972 -1608
rect 2466 -1820 2522 -1384
rect 3559 -1441 3589 -802
rect 3773 -962 3823 833
rect 3896 832 3906 833
rect 3986 832 3996 900
rect 4270 844 4280 898
rect 4340 844 4350 898
rect 4460 846 4470 900
rect 4530 846 4540 900
rect 4722 784 4770 1260
rect 5234 1256 5280 1718
rect 7802 1710 9149 1840
rect 5932 1564 5942 1676
rect 6094 1564 6104 1676
rect 8949 1675 9149 1710
rect 6878 1618 8180 1624
rect 6004 1348 6044 1564
rect 6878 1554 6890 1618
rect 8168 1554 8180 1618
rect 6878 1548 8180 1554
rect 6898 1486 8164 1548
rect 5512 1308 6044 1348
rect 5480 1256 5490 1262
rect 5234 1210 5490 1256
rect 5480 1208 5490 1210
rect 5550 1208 5560 1262
rect 5670 1210 5680 1264
rect 5740 1210 5750 1264
rect 5188 872 5198 950
rect 5270 872 5280 950
rect 5576 898 5586 952
rect 5646 898 5656 952
rect 5766 898 5776 952
rect 5836 898 5846 952
rect 4184 736 4770 784
rect 4152 690 4558 696
rect 4152 644 4164 690
rect 4546 662 4558 690
rect 4546 644 4562 662
rect 4152 638 4562 644
rect 4162 602 4562 638
rect 4174 598 4562 602
rect 4174 568 4552 598
rect 4174 484 4542 568
rect 4182 476 4542 484
rect 4182 454 4304 476
rect 4294 400 4304 454
rect 4386 454 4542 476
rect 4386 400 4396 454
rect 5213 31 5263 872
rect 6004 838 6044 1308
rect 5520 798 6044 838
rect 5466 742 5872 748
rect 5466 696 5478 742
rect 5860 696 5872 742
rect 5466 690 5872 696
rect 5478 656 5860 690
rect 5484 599 5854 656
rect 7350 599 7500 1486
rect 5484 586 7500 599
rect 5504 541 7500 586
rect 5504 500 7450 541
rect 5504 484 5620 500
rect 5610 424 5620 484
rect 5702 484 7450 500
rect 5702 424 5712 484
rect 5213 -19 5575 31
rect 5340 -422 5350 -356
rect 5422 -422 5432 -356
rect 5362 -870 5406 -422
rect 4004 -914 5416 -870
rect 3980 -962 3990 -960
rect 3770 -1012 3990 -962
rect 3980 -1014 3990 -1012
rect 4050 -1014 4060 -960
rect 4174 -1014 4184 -960
rect 4244 -1014 4254 -960
rect 4366 -1016 4376 -962
rect 4436 -1016 4446 -962
rect 4556 -1014 4566 -960
rect 4626 -1014 4636 -960
rect 4748 -1012 4758 -958
rect 4818 -1012 4828 -958
rect 4942 -1012 4952 -958
rect 5012 -1012 5022 -958
rect 5134 -1010 5144 -956
rect 5204 -1010 5214 -956
rect 2789 -1471 3589 -1441
rect 3734 -1510 3744 -1420
rect 3834 -1510 3844 -1420
rect 4076 -1492 4086 -1438
rect 4146 -1492 4156 -1438
rect 4270 -1488 4280 -1434
rect 4340 -1488 4350 -1434
rect 4460 -1484 4470 -1430
rect 4530 -1484 4540 -1430
rect 4654 -1482 4664 -1428
rect 4724 -1482 4734 -1428
rect 4846 -1480 4856 -1426
rect 4916 -1480 4926 -1426
rect 5036 -1478 5046 -1424
rect 5106 -1478 5116 -1424
rect 2730 -1516 3426 -1510
rect 2730 -1568 2742 -1516
rect 3414 -1568 3426 -1516
rect 2730 -1574 3426 -1568
rect 2760 -1820 3384 -1574
rect 3744 -1820 3800 -1510
rect 5364 -1550 5408 -914
rect 5525 -942 5575 -19
rect 8324 -424 8334 -358
rect 8406 -424 8416 -358
rect 8345 -856 8395 -424
rect 5876 -906 8400 -856
rect 5764 -942 5774 -940
rect 5525 -992 5774 -942
rect 5764 -994 5774 -992
rect 5834 -994 5844 -940
rect 5956 -992 5966 -938
rect 6026 -992 6036 -938
rect 6152 -994 6162 -940
rect 6222 -994 6232 -940
rect 6342 -994 6352 -940
rect 6412 -994 6422 -940
rect 6534 -992 6544 -938
rect 6604 -992 6614 -938
rect 6726 -994 6736 -940
rect 6796 -994 6806 -940
rect 6918 -994 6928 -940
rect 6988 -994 6998 -940
rect 7110 -994 7120 -940
rect 7180 -994 7190 -940
rect 7302 -994 7312 -940
rect 7372 -994 7382 -940
rect 7492 -994 7502 -940
rect 7562 -994 7572 -940
rect 7684 -994 7694 -940
rect 7754 -994 7764 -940
rect 7876 -994 7886 -940
rect 7946 -994 7956 -940
rect 8070 -994 8080 -940
rect 8140 -994 8150 -940
rect 5520 -1522 5530 -1432
rect 5620 -1522 5630 -1432
rect 5860 -1496 5870 -1442
rect 5930 -1496 5940 -1442
rect 6052 -1496 6062 -1442
rect 6122 -1496 6132 -1442
rect 6244 -1502 6254 -1448
rect 6314 -1502 6324 -1448
rect 6436 -1498 6446 -1444
rect 6506 -1498 6516 -1444
rect 6628 -1496 6638 -1442
rect 6698 -1496 6708 -1442
rect 6822 -1498 6832 -1444
rect 6892 -1498 6902 -1444
rect 7014 -1500 7024 -1446
rect 7084 -1500 7094 -1446
rect 7206 -1498 7216 -1444
rect 7276 -1498 7286 -1444
rect 7396 -1500 7406 -1446
rect 7466 -1500 7476 -1446
rect 7588 -1502 7598 -1448
rect 7658 -1502 7668 -1448
rect 7780 -1504 7790 -1450
rect 7850 -1504 7860 -1450
rect 7972 -1502 7982 -1448
rect 8042 -1502 8052 -1448
rect 3980 -1594 5408 -1550
rect 3966 -1634 5232 -1628
rect 3966 -1686 3978 -1634
rect 5220 -1686 5232 -1634
rect 3966 -1692 5232 -1686
rect 3974 -1820 5208 -1692
rect 5546 -1784 5602 -1522
rect 8343 -1571 8393 -906
rect 5787 -1621 8393 -1571
rect 5748 -1666 8172 -1660
rect 5748 -1720 5760 -1666
rect 8160 -1720 8172 -1666
rect 5748 -1726 8172 -1720
rect 5768 -1784 8104 -1726
rect 5546 -1820 8104 -1784
rect -106 -1824 8104 -1820
rect -106 -1876 8046 -1824
rect -54 -1996 8046 -1876
rect -54 -2084 5874 -1996
rect -54 -2102 2970 -2084
rect 2742 -2574 2970 -2102
<< via1 >>
rect 2092 1916 2288 2048
rect 3378 1856 3498 1936
rect 4676 1836 4796 1916
rect 5958 1866 6078 1946
rect 2068 1546 2294 1674
rect 1648 1084 1700 1144
rect 1846 1082 1898 1142
rect 992 -488 1152 -302
rect 154 -922 214 -868
rect 348 -916 408 -862
rect -104 -1374 -40 -1304
rect 250 -1366 310 -1312
rect 444 -1362 504 -1308
rect 792 -878 898 -780
rect 1400 832 1466 902
rect 1750 828 1802 888
rect 1942 834 1994 894
rect 3376 1554 3504 1660
rect 2844 1128 2904 1182
rect 3042 1132 3102 1186
rect 2556 848 2630 908
rect 2946 852 3006 906
rect 3138 850 3198 904
rect 1774 410 1850 486
rect 2178 -424 2250 -358
rect 1630 -956 1690 -902
rect 1824 -954 1884 -900
rect 1352 -1422 1442 -1332
rect 1726 -1396 1786 -1342
rect 1920 -1394 1980 -1340
rect 4678 1586 4802 1674
rect 4180 1152 4240 1206
rect 4374 1154 4434 1208
rect 2990 398 3066 474
rect 3540 -426 3612 -360
rect 2752 -918 2812 -864
rect 2948 -916 3008 -862
rect 3140 -912 3200 -858
rect 3332 -912 3392 -858
rect 2462 -1384 2552 -1294
rect 2852 -1362 2912 -1308
rect 3044 -1360 3104 -1306
rect 3238 -1354 3298 -1300
rect 3906 832 3986 900
rect 4280 844 4340 898
rect 4470 846 4530 900
rect 5942 1564 6094 1676
rect 5490 1208 5550 1262
rect 5680 1210 5740 1264
rect 5198 872 5270 950
rect 5586 898 5646 952
rect 5776 898 5836 952
rect 4304 400 4386 476
rect 5620 424 5702 500
rect 5350 -422 5422 -356
rect 3990 -1014 4050 -960
rect 4184 -1014 4244 -960
rect 4376 -1016 4436 -962
rect 4566 -1014 4626 -960
rect 4758 -1012 4818 -958
rect 4952 -1012 5012 -958
rect 5144 -1010 5204 -956
rect 3744 -1510 3834 -1420
rect 4086 -1492 4146 -1438
rect 4280 -1488 4340 -1434
rect 4470 -1484 4530 -1430
rect 4664 -1482 4724 -1428
rect 4856 -1480 4916 -1426
rect 5046 -1478 5106 -1424
rect 8334 -424 8406 -358
rect 5774 -994 5834 -940
rect 5966 -992 6026 -938
rect 6162 -994 6222 -940
rect 6352 -994 6412 -940
rect 6544 -992 6604 -938
rect 6736 -994 6796 -940
rect 6928 -994 6988 -940
rect 7120 -994 7180 -940
rect 7312 -994 7372 -940
rect 7502 -994 7562 -940
rect 7694 -994 7754 -940
rect 7886 -994 7946 -940
rect 8080 -994 8140 -940
rect 5530 -1522 5620 -1432
rect 5870 -1496 5930 -1442
rect 6062 -1496 6122 -1442
rect 6254 -1502 6314 -1448
rect 6446 -1498 6506 -1444
rect 6638 -1496 6698 -1442
rect 6832 -1498 6892 -1444
rect 7024 -1500 7084 -1446
rect 7216 -1498 7276 -1444
rect 7406 -1500 7466 -1446
rect 7598 -1502 7658 -1448
rect 7790 -1504 7850 -1450
rect 7982 -1502 8042 -1448
<< metal2 >>
rect 2092 2048 2288 2056
rect 5958 1946 6078 1956
rect 2092 1906 2288 1916
rect 3378 1936 3498 1946
rect 2136 1684 2242 1906
rect 3378 1846 3498 1856
rect 4676 1916 4796 1926
rect 2068 1674 2294 1684
rect 3400 1670 3474 1846
rect 5958 1856 6078 1866
rect 4676 1826 4796 1836
rect 4708 1684 4782 1826
rect 5980 1686 6048 1856
rect 4678 1674 4802 1684
rect 2068 1536 2294 1546
rect 3376 1660 3504 1670
rect 4678 1576 4802 1586
rect 5942 1676 6094 1686
rect 5942 1554 6094 1564
rect 3376 1544 3504 1554
rect 5490 1262 5550 1272
rect 4180 1206 4240 1216
rect 2844 1182 2904 1192
rect 1648 1144 1700 1154
rect 1846 1142 1898 1152
rect 1700 1094 1846 1132
rect 1648 1074 1700 1084
rect 3042 1186 3102 1196
rect 2904 1144 3042 1174
rect 2844 1118 2904 1128
rect 4374 1208 4434 1218
rect 4240 1158 4374 1194
rect 4180 1142 4240 1152
rect 5680 1264 5740 1274
rect 5550 1216 5680 1256
rect 5490 1198 5550 1208
rect 5680 1200 5740 1210
rect 4374 1144 4434 1154
rect 3042 1122 3102 1132
rect 1846 1072 1898 1082
rect 5198 950 5270 960
rect 1400 902 1466 912
rect 2556 908 2630 918
rect 1750 888 1802 898
rect 1466 846 1750 880
rect 1400 822 1466 832
rect 1942 894 1994 904
rect 1802 846 1942 880
rect 1750 818 1802 828
rect 2946 906 3006 916
rect 2630 864 2946 894
rect 2556 838 2630 848
rect 3138 904 3198 914
rect 3006 864 3138 894
rect 2946 842 3006 852
rect 3138 840 3198 850
rect 3906 900 3986 910
rect 1942 824 1994 834
rect 4280 898 4340 908
rect 3986 846 4280 888
rect 4470 900 4530 910
rect 4340 846 4470 888
rect 5586 952 5646 962
rect 5270 900 5586 936
rect 5776 952 5836 962
rect 5646 900 5776 936
rect 5586 888 5646 898
rect 5776 888 5836 898
rect 5198 862 5270 872
rect 4280 834 4340 844
rect 4470 836 4530 846
rect 3906 822 3986 832
rect 5620 500 5702 510
rect 1774 486 1850 496
rect 808 440 884 442
rect 808 410 1774 440
rect 2990 474 3066 484
rect 1850 410 2990 440
rect 808 398 2990 410
rect 4304 476 4386 486
rect 3066 400 4304 440
rect 4386 424 5620 440
rect 5702 424 5772 440
rect 4386 400 5772 424
rect 3066 398 5772 400
rect 808 364 5772 398
rect 808 -770 884 364
rect 992 -302 1152 -292
rect 1152 -356 8430 -336
rect 1152 -358 5350 -356
rect 1152 -424 2178 -358
rect 2250 -360 5350 -358
rect 2250 -424 3540 -360
rect 1152 -426 3540 -424
rect 3612 -422 5350 -360
rect 5422 -358 8430 -356
rect 5422 -422 8334 -358
rect 3612 -424 8334 -422
rect 8406 -424 8430 -358
rect 3612 -426 8430 -424
rect 1152 -442 8430 -426
rect 992 -498 1152 -488
rect 792 -780 898 -770
rect 154 -868 214 -858
rect 348 -862 408 -852
rect 214 -910 348 -868
rect 154 -932 214 -922
rect 792 -888 898 -878
rect 2752 -864 2812 -854
rect 348 -926 408 -916
rect 1630 -902 1690 -892
rect 1824 -900 1884 -890
rect 1690 -952 1824 -906
rect 1630 -966 1690 -956
rect 2948 -862 3008 -852
rect 2812 -912 2948 -866
rect 2752 -928 2812 -918
rect 3140 -858 3200 -848
rect 3008 -912 3140 -866
rect 3332 -858 3392 -848
rect 3200 -912 3332 -866
rect 2948 -926 3008 -916
rect 3140 -922 3200 -912
rect 3332 -922 3392 -912
rect 5774 -940 5834 -930
rect 1824 -964 1884 -954
rect 3990 -960 4050 -950
rect 3962 -1008 3990 -966
rect 4184 -960 4244 -950
rect 4050 -1008 4184 -966
rect 3990 -1024 4050 -1014
rect 4376 -962 4436 -952
rect 4244 -1008 4376 -966
rect 4184 -1024 4244 -1014
rect 4566 -960 4626 -950
rect 4436 -1008 4566 -966
rect 4376 -1026 4436 -1016
rect 4758 -958 4818 -948
rect 4626 -1008 4758 -966
rect 4566 -1024 4626 -1014
rect 4952 -958 5012 -948
rect 4818 -1008 4952 -966
rect 4758 -1022 4818 -1012
rect 5144 -956 5204 -946
rect 5012 -1008 5144 -966
rect 4952 -1022 5012 -1012
rect 5740 -988 5774 -946
rect 5966 -938 6026 -928
rect 5834 -988 5966 -946
rect 5774 -1004 5834 -994
rect 6162 -940 6222 -930
rect 6026 -988 6162 -946
rect 5966 -1002 6026 -992
rect 6352 -940 6412 -930
rect 6222 -988 6352 -946
rect 6162 -1004 6222 -994
rect 6544 -938 6604 -928
rect 6412 -988 6544 -946
rect 6352 -1004 6412 -994
rect 6736 -940 6796 -930
rect 6604 -988 6736 -946
rect 6544 -1002 6604 -992
rect 6928 -940 6988 -930
rect 6796 -988 6928 -946
rect 6736 -1004 6796 -994
rect 7120 -940 7180 -930
rect 6988 -988 7120 -946
rect 6928 -1004 6988 -994
rect 7312 -940 7372 -930
rect 7180 -988 7312 -946
rect 7120 -1004 7180 -994
rect 7502 -940 7562 -930
rect 7372 -988 7502 -946
rect 7312 -1004 7372 -994
rect 7694 -940 7754 -930
rect 7562 -988 7694 -946
rect 7502 -1004 7562 -994
rect 7886 -940 7946 -930
rect 7754 -988 7886 -946
rect 7694 -1004 7754 -994
rect 8080 -940 8140 -930
rect 7946 -988 8080 -946
rect 7886 -1004 7946 -994
rect 8080 -1004 8140 -994
rect 5144 -1020 5204 -1010
rect 2462 -1294 2552 -1284
rect -104 -1304 -40 -1294
rect 250 -1312 310 -1302
rect -40 -1362 250 -1318
rect -104 -1384 -40 -1374
rect 444 -1308 504 -1298
rect 310 -1362 444 -1318
rect 250 -1376 310 -1366
rect 444 -1372 504 -1362
rect 1352 -1332 1442 -1322
rect 1726 -1342 1786 -1332
rect 1442 -1396 1726 -1354
rect 1920 -1340 1980 -1330
rect 1786 -1394 1920 -1354
rect 2852 -1308 2912 -1298
rect 2552 -1358 2852 -1316
rect 3044 -1306 3104 -1296
rect 2912 -1358 3044 -1316
rect 2852 -1372 2912 -1362
rect 3238 -1300 3298 -1290
rect 3104 -1354 3238 -1316
rect 3104 -1358 3298 -1354
rect 3044 -1370 3104 -1360
rect 3238 -1364 3298 -1358
rect 2462 -1394 2552 -1384
rect 1786 -1396 1980 -1394
rect 1442 -1400 1980 -1396
rect 1726 -1406 1786 -1400
rect 1920 -1404 1980 -1400
rect 1352 -1432 1442 -1422
rect 3744 -1420 3834 -1410
rect 4086 -1436 4146 -1428
rect 4280 -1434 4340 -1424
rect 3834 -1438 4280 -1436
rect 3834 -1484 4086 -1438
rect 4146 -1484 4280 -1438
rect 4086 -1502 4146 -1492
rect 4470 -1430 4530 -1420
rect 4340 -1484 4470 -1436
rect 4664 -1428 4724 -1418
rect 4530 -1482 4664 -1436
rect 4856 -1426 4916 -1416
rect 4724 -1480 4856 -1436
rect 5046 -1424 5106 -1414
rect 4916 -1478 5046 -1436
rect 4916 -1480 5106 -1478
rect 4724 -1482 5106 -1480
rect 4530 -1484 5106 -1482
rect 4280 -1498 4340 -1488
rect 4470 -1494 4530 -1484
rect 4664 -1492 4724 -1484
rect 4856 -1490 4916 -1484
rect 5046 -1488 5106 -1484
rect 5530 -1432 5620 -1422
rect 3744 -1520 3834 -1510
rect 5870 -1442 5930 -1432
rect 5620 -1496 5870 -1458
rect 6062 -1442 6122 -1432
rect 5930 -1496 6062 -1458
rect 6254 -1448 6314 -1438
rect 6122 -1496 6254 -1458
rect 5870 -1506 5930 -1496
rect 6062 -1506 6122 -1496
rect 6446 -1444 6506 -1434
rect 6314 -1496 6446 -1458
rect 6254 -1512 6314 -1502
rect 6638 -1442 6698 -1432
rect 6506 -1496 6638 -1458
rect 6832 -1444 6892 -1434
rect 6698 -1496 6832 -1458
rect 6446 -1508 6506 -1498
rect 6638 -1506 6698 -1496
rect 7024 -1446 7084 -1436
rect 6892 -1496 7024 -1458
rect 6832 -1508 6892 -1498
rect 7216 -1444 7276 -1434
rect 7084 -1496 7216 -1458
rect 7024 -1510 7084 -1500
rect 7406 -1446 7466 -1436
rect 7276 -1496 7406 -1458
rect 7216 -1508 7276 -1498
rect 7598 -1448 7658 -1438
rect 7466 -1496 7598 -1458
rect 7406 -1510 7466 -1500
rect 7790 -1450 7850 -1440
rect 7658 -1496 7790 -1458
rect 7598 -1512 7658 -1502
rect 7982 -1448 8042 -1438
rect 7850 -1496 7982 -1458
rect 7790 -1514 7850 -1504
rect 7982 -1512 8042 -1502
rect 5530 -1532 5620 -1522
use sky130_fd_pr__nfet_01v8_lvt_HMT3AU  XN1
timestamp 1751989567
transform 1 0 1823 0 1 1018
box -311 -410 311 410
use sky130_fd_pr__nfet_01v8_lvt_HMT3AU  XN2
timestamp 1751989567
transform 1 0 3023 0 1 1032
box -311 -410 311 410
use sky130_fd_pr__nfet_01v8_lvt_HMT3AU  XN3
timestamp 1751989567
transform 1 0 4355 0 1 1024
box -311 -410 311 410
use sky130_fd_pr__nfet_01v8_lvt_HMT3AU  XN4
timestamp 1751989567
transform 1 0 5663 0 1 1076
box -311 -410 311 410
use sky130_fd_pr__nfet_01v8_lvt_HFZZWY  XQ0
timestamp 1751989567
transform 1 0 329 0 1 -1123
box -311 -477 311 477
use sky130_fd_pr__nfet_01v8_lvt_HFZZWY  XQ1
timestamp 1751989567
transform 1 0 1805 0 1 -1151
box -311 -477 311 477
use sky130_fd_pr__nfet_01v8_lvt_EEV8MN  XQ2
timestamp 1751989567
transform 1 0 3073 0 1 -1115
box -455 -477 455 477
use sky130_fd_pr__nfet_01v8_lvt_34GFY5  XQ3
timestamp 1751989567
transform 1 0 4597 0 1 -1227
box -743 -485 743 485
use sky130_fd_pr__nfet_01v8_lvt_GYBLDK  XQ4
timestamp 1751989567
transform 1 0 6957 0 1 -1222
box -1319 -498 1319 498
use sky130_fd_pr__res_xhigh_po_0p35_48NHYL  XR3
timestamp 1751989567
transform 1 0 -1739 0 1 970
box -201 -2182 201 2182
use sky130_fd_pr__res_xhigh_po_0p35_48NHYL  XR4
timestamp 1751989567
transform 1 0 -1151 0 1 970
box -201 -2182 201 2182
use sky130_fd_pr__res_xhigh_po_0p69_NP4GWP  XR5
timestamp 1751989567
transform 0 -1 7525 1 0 1773
box -235 -757 235 757
<< labels >>
flabel metal1 6412 1836 6612 2036 0 FreeSans 256 0 0 0 OUT
port 5 nsew
flabel metal1 8949 1675 9149 1875 0 FreeSans 256 0 0 0 VDD
port 6 nsew
flabel metal1 -2462 -942 -2262 -742 0 FreeSans 256 0 0 0 Vref
port 4 nsew
flabel metal1 2088 2124 2288 2324 0 FreeSans 256 0 0 0 D0
port 2 nsew
flabel metal1 3334 2044 3534 2244 0 FreeSans 256 0 0 0 D1
port 3 nsew
flabel metal1 4618 1972 4818 2172 0 FreeSans 256 0 0 0 D2
port 1 nsew
flabel metal1 5914 2012 6114 2212 0 FreeSans 256 0 0 0 D3
port 0 nsew
flabel metal1 2742 -2574 2970 -2298 0 FreeSans 480 0 0 0 VSS
port 9 nsew
<< end >>
